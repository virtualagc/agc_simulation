`timescale 1ns/1ps
`default_nettype none

module fpga_ch77_alarm_box(p4VDC, p4VSW, GND, SIM_RST, SIM_CLK, MCTRAL_n, MPAL_n, MRCH, MRPTAL_n, MSCAFL_n, MSCDBL_n, MT01, MT05, MT12, MTCAL_n, MVFAIL_n, MWATCH_n, MWCH, MWL01, MWL02, MWL03, MWL04, MWL05, MWL06, MWSG, DBLTST, DOSCAL, MAMU, MDT01, MDT02, MDT03, MDT04, MDT05, MDT06, MDT07, MDT08, MDT09, MDT10, MDT11, MDT12, MDT13, MDT14, MDT15, MDT16, MLDCH, MLOAD, MNHNC, MNHRPT, MNHSBF, MONPAR, MONWBK, MRDCH, MREAD, MSBSTP, MSTP, MSTRT, MTCSAI, NHALGA);
    input wire p4VDC;
    input wire p4VSW;
    input wire GND;
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire MCTRAL_n;
    input wire MPAL_n;
    input wire MRCH;
    input wire MRPTAL_n;
    input wire MSCAFL_n;
    input wire MSCDBL_n;
    input wire MT01;
    input wire MT05;
    input wire MT12;
    input wire MTCAL_n;
    input wire MVFAIL_n;
    input wire MWATCH_n;
    input wire MWCH;
    input wire MWL01;
    input wire MWL02;
    input wire MWL03;
    input wire MWL04;
    input wire MWL05;
    input wire MWL06;
    input wire MWSG;
    output wire DBLTST;
    output wire DOSCAL;
    output wire MAMU;
    output wire MDT01;
    output wire MDT02;
    output wire MDT03;
    output wire MDT04;
    output wire MDT05;
    output wire MDT06;
    output wire MDT07;
    output wire MDT08;
    output wire MDT09;
    output wire MDT10;
    output wire MDT11;
    output wire MDT12;
    output wire MDT13;
    output wire MDT14;
    output wire MDT15;
    output wire MDT16;
    output wire MLDCH;
    output wire MLOAD;
    output wire MNHNC;
    output wire MNHRPT;
    output wire MNHSBF;
    output wire MONPAR;
    output wire MONWBK;
    output wire MRDCH;
    output wire MREAD;
    output wire MSBSTP;
    output wire MSTP;
    output wire MSTRT;
    output wire MTCSAI;
    output wire NHALGA;
    wire __RestartMonitor__CCH77;
    wire __RestartMonitor__RCH77_n;
    wand __Z99_NET_100;
    wire __Z99_NET_100_U77004_2;
    wire __Z99_NET_100_U77004_4;
    wire __Z99_NET_101;
    wire __Z99_NET_102;
    wire __Z99_NET_105;
    wire __Z99_NET_56;
    wire __Z99_NET_57;
    wire __Z99_NET_58;
    wire __Z99_NET_59;
    wire __Z99_NET_60;
    wire __Z99_NET_61;
    wire __Z99_NET_62;
    wire __Z99_NET_63;
    wire __Z99_NET_64;
    wire __Z99_NET_65;
    wire __Z99_NET_66;
    wire __Z99_NET_67;
    wire __Z99_NET_68;
    wire __Z99_NET_69;
    wire __Z99_NET_70;
    wire __Z99_NET_71;
    wire __Z99_NET_72;
    wire __Z99_NET_73;
    wire __Z99_NET_74;
    wire __Z99_NET_75;
    wire __Z99_NET_76;
    wire __Z99_NET_77;
    wire __Z99_NET_78;
    wire __Z99_NET_79;
    wire __Z99_NET_80;
    wire __Z99_NET_81;
    wire __Z99_NET_82;
    wire __Z99_NET_83;
    wire __Z99_NET_84;
    wire __Z99_NET_87;
    wire __Z99_NET_88;
    wire __Z99_NET_89;
    wire __Z99_NET_90;
    wire __Z99_NET_91;
    wire __Z99_NET_92;
    wire __Z99_NET_94;
    wire __Z99_NET_95;
    wire __Z99_NET_96;
    wire __Z99_NET_98;
    wire __Z99_NET_99;

    assign MDT10 = GND;
    assign MDT11 = GND;
    assign MDT12 = GND;
    assign MDT13 = GND;
    assign MDT14 = GND;
    assign MDT15 = GND;
    assign MDT16 = GND;
    assign MNHSBF = GND;
    assign MNHNC = GND;
    assign MNHRPT = GND;
    assign MTCSAI = GND;
    assign MSTRT = GND;
    assign MSTP = GND;
    assign MSBSTP = GND;
    assign MRDCH = GND;
    assign MLDCH = GND;
    assign MONPAR = GND;
    assign MONWBK = GND;
    assign MLOAD = GND;
    assign MREAD = GND;
    assign NHALGA = GND;
    assign DOSCAL = GND;
    assign DBLTST = GND;
    assign MAMU = GND;
    U74HC04 U77001(MWL01, __Z99_NET_102, MWL02, __Z99_NET_91, MWL03, __Z99_NET_92, GND, __Z99_NET_105, MWL04, __Z99_NET_89, MWL05, __Z99_NET_90, MWL06, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0) U77002(MT01, __Z99_NET_101, MWSG, __Z99_NET_94, MWCH, __Z99_NET_87, GND, __Z99_NET_88, MRCH, __RestartMonitor__RCH77_n, __Z99_NET_73, __Z99_NET_75, MPAL_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U77003(__Z99_NET_96, __Z99_NET_102, __Z99_NET_91, __Z99_NET_92, __Z99_NET_105,  , GND,  , __Z99_NET_89, __Z99_NET_90, __Z99_NET_101, __Z99_NET_94, __Z99_NET_95, p4VSW, SIM_RST, SIM_CLK);
    assign __Z99_NET_100 = __Z99_NET_100_U77004_2;
    assign __Z99_NET_100 = __Z99_NET_100_U77004_4;
    U74LVC07 U77004(__Z99_NET_96, __Z99_NET_100_U77004_2, __Z99_NET_95, __Z99_NET_100_U77004_4,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U77005(__Z99_NET_98, MT12, __Z99_NET_99, __Z99_NET_99, __Z99_NET_98, __Z99_NET_100, GND, __Z99_NET_88, __Z99_NET_99, __Z99_NET_73, __Z99_NET_87, __Z99_NET_99, __RestartMonitor__CCH77, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U77006(__Z99_NET_56, __Z99_NET_75, __Z99_NET_74, __Z99_NET_74, __Z99_NET_56, __RestartMonitor__CCH77, GND, __Z99_NET_69, __Z99_NET_76, __Z99_NET_64, __Z99_NET_64, __RestartMonitor__CCH77, __Z99_NET_76, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U77007(__Z99_NET_69, MPAL_n, __Z99_NET_70, __Z99_NET_65, __Z99_NET_72, __Z99_NET_71, GND, __Z99_NET_65, __RestartMonitor__CCH77, __Z99_NET_71, __Z99_NET_82, __Z99_NET_81, __Z99_NET_66, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U77008(MT05, __Z99_NET_70, MTCAL_n, __Z99_NET_72, MRPTAL_n, __Z99_NET_82, GND, __Z99_NET_84, MWATCH_n, __Z99_NET_78, MVFAIL_n, __Z99_NET_80, MCTRAL_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U77009(__Z99_NET_81, __Z99_NET_66, __RestartMonitor__CCH77, __Z99_NET_63, __Z99_NET_84, __Z99_NET_83, GND, __Z99_NET_63, __RestartMonitor__CCH77, __Z99_NET_83, __Z99_NET_78, __Z99_NET_77, __Z99_NET_67, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U77010(__Z99_NET_77, __Z99_NET_67, __RestartMonitor__CCH77, __Z99_NET_68, __Z99_NET_80, __Z99_NET_79, GND, __Z99_NET_68, __RestartMonitor__CCH77, __Z99_NET_79, __Z99_NET_59, __Z99_NET_57, __Z99_NET_58, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U77011(__Z99_NET_57, __Z99_NET_58, __RestartMonitor__CCH77, __Z99_NET_62, __Z99_NET_60, __Z99_NET_61, GND, __Z99_NET_62, __RestartMonitor__CCH77, __Z99_NET_61,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U77012(MSCAFL_n, __Z99_NET_59, MSCDBL_n, __Z99_NET_60,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U77013(__RestartMonitor__RCH77_n, __Z99_NET_56, __RestartMonitor__RCH77_n, __Z99_NET_64, GND, MDT02, GND, MDT03, __RestartMonitor__RCH77_n, __Z99_NET_65, GND, MDT01, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U77014(__RestartMonitor__RCH77_n, __Z99_NET_66, __RestartMonitor__RCH77_n, __Z99_NET_63, GND, MDT05, GND, MDT06, __RestartMonitor__RCH77_n, __Z99_NET_67, GND, MDT04, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U77015(__RestartMonitor__RCH77_n, __Z99_NET_68, __RestartMonitor__RCH77_n, __Z99_NET_58, GND, MDT08, GND, MDT09, __RestartMonitor__RCH77_n, __Z99_NET_62, GND, MDT07, GND, p4VSW, SIM_RST, SIM_CLK);
endmodule
