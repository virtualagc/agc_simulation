`timescale 1ns/1ps

module stage_branch(VCC, GND, SIM_RST, GOJAM, PHS2_n, PHS3_n, PHS4, PHS4_n, T01, T03, T01_n, T02_n, T03_n, T04_n, T05_n, T06_n, T07_n, T08_n, T09_n, T10_n, T11_n, T12_n, SQ0_n, SQ1_n, SQ2_n, QC0_n, QC1_n, QC2_n, QC3_n, SQEXT_n, SQR10, SQR10_n, SQR12_n, STRTFC, WL16_n, WL15_n, WL14_n, WL13_n, WL12_n, WL11_n, WL10_n, WL09_n, WL08_n, WL07_n, WL06_n, WL05_n, WL04_n, WL03_n, WL02_n, WL01_n, OVF_n, UNF_n, SUMA16_n, SUMB16_n, EXST0_n, EXST1_n, ST1, ST2, RSTSTG, TMZ_n, TOV_n, TSGN_n, TSGU_n, TPZG_n, DVST, GEQZRO_n, TRSM, NDR100_n, INKL, L15_n, TL15, XT1_n, XB7_n, MTCSAI, MP0_n, MP1, MP3A, MP3_n, IC12, IC13, IC15, TS0_n, RSM3, RSM3_n, STORE1_n, n7XP14, ST0_n, ST1_n, STD2, ST3_n, ST4_n, BR2_n, BR1B2B, KRPT, RXOR0, n5XP4);
    input wire SIM_RST;
    output wire BR1B2B;
    output wire BR2_n;
    input wire DVST;
    input wire EXST0_n;
    input wire EXST1_n;
    input wire GEQZRO_n;
    input wire GND;
    input wire GOJAM;
    input wire IC12;
    input wire IC13;
    input wire IC15;
    input wire INKL;
    output wire KRPT;
    input wire L15_n;
    input wire MP0_n;
    input wire MP1;
    input wire MP3A;
    input wire MP3_n;
    input wire MTCSAI;
    input wire NDR100_n;
    wire NET_182;
    wire NET_183;
    wire NET_184;
    wire NET_185;
    wire NET_186;
    wire NET_187;
    wire NET_188;
    wire NET_189;
    wire NET_190;
    wire NET_191;
    wire NET_192;
    wire NET_193;
    wire NET_194;
    wire NET_195;
    wire NET_196;
    wire NET_197;
    wire NET_198;
    wire NET_199;
    wire NET_200;
    wire NET_201;
    wire NET_202;
    wire NET_203;
    wire NET_204;
    wire NET_205;
    wire NET_206;
    wire NET_207;
    wire NET_210;
    wire NET_211;
    wire NET_214;
    wire NET_215;
    wire NET_216;
    wire NET_217;
    wire NET_218;
    wire NET_219;
    wire NET_220;
    wire NET_221;
    wire NET_224;
    wire NET_225;
    wire NET_226;
    wire NET_227;
    wire NET_228;
    wire NET_229;
    wire NET_230;
    wire NET_231;
    wire NET_232;
    wire NET_233;
    wire NET_234;
    wire NET_235;
    wire NET_236;
    wire NET_237;
    wire NET_238;
    wire NET_239;
    wire NET_240;
    wire NET_241;
    wire NET_242;
    wire NET_243;
    wire NET_244;
    wire NET_245;
    wire NET_246;
    wire NET_247;
    wire NET_248;
    wire NET_249;
    wire NET_250;
    wire NET_251;
    wire NET_252;
    wire NET_253;
    wire NET_254;
    wire NET_255;
    wire NET_258;
    wire NET_259;
    wire NET_260;
    wire NET_261;
    wire NET_262;
    wire NET_263;
    wire NET_264;
    wire NET_265;
    wire NET_266;
    wire NET_267;
    wire NET_268;
    wire NET_269;
    wire NET_271;
    wire NET_272;
    wire NET_273;
    wire NET_274;
    wire NET_275;
    wire NET_276;
    wire NET_277;
    wire NET_278;
    wire NET_279;
    wire NET_280;
    wire NET_281;
    wire NET_282;
    wire NET_283;
    wire NET_284;
    wire NET_285;
    wire NET_286;
    wire NET_287;
    wire NET_288;
    wire NET_289;
    wire NET_290;
    wire NET_291;
    wire NET_292;
    wire NET_293;
    wire NET_294;
    wire NET_295;
    wire NET_296;
    wire NET_297;
    wire NET_298;
    wire NET_299;
    wire NET_300;
    wire NET_301;
    wire NET_302;
    wire NET_303;
    wire NET_304;
    wire NET_305;
    wire NET_306;
    wire NET_307;
    wire NET_308;
    wire NET_309;
    wire NET_310;
    wire NET_311;
    wire NET_312;
    wire NET_313;
    wire NET_314;
    wire NET_315;
    wire NET_316;
    wire NET_317;
    wire NET_318;
    wire NET_319;
    wire NET_320;
    wire NET_321;
    wire NET_322;
    wire NET_323;
    wire NET_324;
    wire NET_327;
    wire NET_328;
    wire NET_329;
    wire NET_330;
    input wire OVF_n;
    input wire PHS2_n;
    input wire PHS3_n;
    input wire PHS4;
    input wire PHS4_n;
    input wire QC0_n;
    input wire QC1_n;
    input wire QC2_n;
    input wire QC3_n;
    input wire RSM3;
    input wire RSM3_n;
    input wire RSTSTG;
    output wire RXOR0;
    input wire SQ0_n;
    input wire SQ1_n;
    input wire SQ2_n;
    input wire SQEXT_n;
    input wire SQR10;
    input wire SQR10_n;
    input wire SQR12_n;
    output wire ST0_n;
    input wire ST1;
    output wire ST1_n;
    input wire ST2;
    output wire ST3_n;
    output wire ST4_n;
    output wire STD2;
    input wire STORE1_n;
    input wire STRTFC;
    input wire SUMA16_n;
    input wire SUMB16_n;
    input wire T01;
    input wire T01_n;
    input wire T02_n;
    input wire T03;
    input wire T03_n;
    input wire T04_n;
    input wire T05_n;
    input wire T06_n;
    input wire T07_n;
    input wire T08_n;
    input wire T09_n;
    input wire T10_n;
    input wire T11_n;
    input wire T12_n;
    output wire TL15;
    inout wire TMZ_n;
    input wire TOV_n;
    input wire TPZG_n;
    input wire TRSM;
    input wire TS0_n;
    inout wire TSGN_n;
    input wire TSGU_n;
    input wire UNF_n;
    input wire VCC;
    input wire WL01_n;
    input wire WL02_n;
    input wire WL03_n;
    input wire WL04_n;
    input wire WL05_n;
    input wire WL06_n;
    input wire WL07_n;
    input wire WL08_n;
    input wire WL09_n;
    input wire WL10_n;
    input wire WL11_n;
    input wire WL12_n;
    input wire WL13_n;
    input wire WL14_n;
    input wire WL15_n;
    input wire WL16_n;
    input wire XB7_n;
    input wire XT1_n;
    wire __A04_1__BR1;
    wire __A04_1__BR1_n;
    wire __A04_1__BR2;
    wire __A04_1__DIVSTG;
    wire __A04_1__DIV_n;
    wire __A04_1__DV0;
    wire __A04_1__DV0_n;
    wire __A04_1__DV1;
    wire __A04_1__DV1376;
    wire __A04_1__DV1736_n;
    wire __A04_1__DV1_n;
    wire __A04_1__DV376;
    wire __A04_1__DV3764;
    wire __A04_1__DV376_n;
    wire __A04_1__DV4;
    wire __A04_1__DV4_n;
    wire __A04_1__MBR1;
    wire __A04_1__MBR2;
    wire __A04_1__MST1;
    wire __A04_1__MST2;
    wire __A04_1__MST3;
    wire __A04_1__SGUM;
    wire __A04_1__ST1376_n;
    wire __A04_1__ST376;
    wire __A04_1__ST376_n;
    wire __A04_1__STG1;
    wire __A04_1__STG2;
    wire __A04_1__STG3;
    wire __A04_1__T12USE_n;
    wire __A04_1__TSGN2;
    wire __A04_2__1XP10;
    wire __A04_2__2XP3;
    wire __A04_2__2XP5;
    wire __A04_2__3XP2;
    wire __A04_2__3XP7;
    wire __A04_2__4XP11;
    wire __A04_2__4XP5;
    wire __A04_2__5XP11;
    wire __A04_2__5XP28;
    wire __A04_2__6XP5;
    wire __A04_2__7XP19;
    wire __A04_2__8PP4;
    wire __A04_2__8XP5;
    wire __A04_2__8XP6;
    wire __A04_2__9XP1;
    wire __A04_2__B15X;
    wire __A04_2__BR12B;
    wire __A04_2__BR12B_n;
    wire __A04_2__BR1B2;
    wire __A04_2__BR1B2B_n;
    wire __A04_2__BR1B2_n;
    wire __A04_2__BRDIF_n;
    wire __A04_2__CI_n;
    wire __A04_2__DV0_n;
    wire __A04_2__INOUT;
    wire __A04_2__INOUT_n;
    wire __A04_2__L16_n;
    wire __A04_2__MP0T10;
    wire __A04_2__MRSC;
    wire __A04_2__PRINC;
    wire __A04_2__R15;
    wire __A04_2__R1C_n;
    wire __A04_2__RAND0;
    wire __A04_2__RA_n;
    wire __A04_2__RB1_n;
    wire __A04_2__RB2;
    wire __A04_2__RB_n;
    wire __A04_2__RC_n;
    wire __A04_2__READ0;
    wire __A04_2__READ0_n;
    wire __A04_2__ROR0;
    wire __A04_2__RRPA;
    wire __A04_2__RSC_n;
    wire __A04_2__RUPT0;
    wire __A04_2__RUPT0_n;
    wire __A04_2__RUPT1;
    wire __A04_2__RUPT1_n;
    wire __A04_2__RXOR0_n;
    wire __A04_2__WAND0;
    wire __A04_2__WCH_n;
    wire __A04_2__WG_n;
    wire __A04_2__WL_n;
    wire __A04_2__WOR0;
    wire __A04_2__WOR0_n;
    wire __A04_2__WRITE0;
    wire __A04_2__WRITE0_n;
    wire __A04_2__WY_n;
    output wire n5XP4;
    input wire n7XP14;

    pullup R3004(NET_215);
    pullup R3005(NET_214);
    pullup R4001(NET_249);
    pullup R4002(NET_237);
    pullup R4003(__A04_1__SGUM);
    pullup R4006(NET_219);
    pullup R4007(NET_207);
    pullup R4008(__A04_2__5XP11);
    pullup R4009(__A04_2__RA_n);
    pullup R4010(__A04_2__WG_n);
    pullup R4011(NET_283);
    pullup R4012(__A04_2__RA_n);
    pullup R4013(TMZ_n);
    pullup R4014(__A04_2__WY_n);
    pullup R4015(__A04_2__WL_n);
    pullup R4016(__A04_2__RC_n);
    pullup R4017(__A04_2__RB_n);
    pullup R4018(__A04_2__CI_n);
    pullup R4019(TSGN_n);
    pullup R4020(__A04_2__RB1_n);
    pullup R4021(__A04_2__L16_n);
    U74HC02 #(0, 0, 0, 1) U4001(__A04_1__T12USE_n, DVST, NET_242, __A04_1__DIVSTG, __A04_1__T12USE_n, T03, GND, NET_243, NET_241, NET_268, GOJAM, MTCSAI, NET_248, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U4002(T03, __A04_1__T12USE_n, __A04_1__T12USE_n, RSTSTG, GOJAM, NET_242, GND, NET_241, PHS3_n, NET_242, T12_n, NET_243, PHS3_n, VCC, SIM_RST);
    U74LVC07 U4003(NET_248, NET_249, NET_247, NET_249, NET_228, NET_237, GND, NET_237, NET_231, __A04_1__SGUM, NET_198, __A04_1__SGUM, NET_197, VCC, SIM_RST);
    U74HC27 #(1, 1, 0) U4004(ST1, NET_244, __A04_1__STG1, __A04_1__STG3, __A04_1__STG2, NET_230, GND, NET_253, __A04_1__STG2, __A04_1__STG3, NET_235, NET_247, NET_246, VCC, SIM_RST);
    U74HC02 U4005(NET_246, NET_249, T01, NET_244, NET_233, NET_264, GND, NET_268, NET_249, NET_240, NET_246, NET_268, NET_245, VCC, SIM_RST);
    U74HC02 #(1, 0, 1, 0) U4006(NET_235, NET_240, __A04_1__STG1, __A04_1__STG1, NET_235, NET_245, GND, ST2, NET_229, NET_228, NET_233, NET_235, NET_234, VCC, SIM_RST);
    U74HC04 U4007(NET_235, __A04_1__MST1, NET_258, __A04_1__MST2, NET_264, __A04_1__MST3, GND, __A04_1__MBR1, NET_215, __A04_1__MBR2, NET_207, NET_233, DVST, VCC, SIM_RST);
    U74HC04 #(0, 1, 1, 1, 0, 0) U4008(NET_230, ST0_n, NET_253, ST1_n, NET_265, ST3_n, GND, ST4_n, NET_251, __A04_1__ST376_n, __A04_1__ST376, __A04_1__DV1736_n, __A04_1__DV1376, VCC, SIM_RST);
    U74HC27 #(1, 0, 0) U4009(NET_234, MTCSAI, NET_237, GOJAM, T01, NET_232, GND, NET_265, __A04_1__STG3, NET_258, NET_235, NET_231, NET_232, VCC, SIM_RST);
    U74HC4002 U4010(NET_229, NET_210, XT1_n, XB7_n, NDR100_n, NET_239, GND, NET_238, NET_255, STRTFC, T01, RSTSTG, NET_260, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U4011(NET_261, NET_268, NET_237, NET_236, NET_232, NET_268, GND, NET_261, __A04_1__STG2, NET_258, NET_258, NET_236, __A04_1__STG2, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U4012(NET_259, NET_233, NET_258, NET_255, NET_259, NET_260, GND, NET_268, NET_255, NET_266, NET_260, NET_268, NET_267, VCC, SIM_RST);
    U74HC02 #(1, 0, 0, 0) U4013(NET_264, NET_266, __A04_1__STG3, __A04_1__STG3, NET_264, NET_267, GND, __A04_1__STG1, __A04_1__STG3, NET_250, NET_258, NET_250, __A04_1__ST376, VCC, SIM_RST);
    U74HC4002 U4014(STD2, INKL, __A04_1__STG1, __A04_1__STG3, NET_258, NET_263, GND, NET_262, SQ0_n, EXST1_n, QC3_n, SQR10_n, __A04_2__RUPT1, VCC, SIM_RST);
    U74HC27 U4015(NET_264, __A04_1__STG1, QC0_n, SQEXT_n, SQ1_n, NET_252, GND, NET_198, SUMB16_n, SUMA16_n, TSGU_n, NET_251, __A04_1__STG2, VCC, SIM_RST);
    U74HC02 U4016(NET_254, NET_251, __A04_1__ST376, __A04_1__DV3764, __A04_1__DIV_n, NET_254, GND, NET_253, __A04_1__ST376, __A04_1__ST1376_n, __A04_1__DIV_n, __A04_1__ST1376_n, __A04_1__DV1376, VCC, SIM_RST);
    U74HC04 U4017(NET_252, __A04_1__DIV_n, __A04_1__DV0, __A04_1__DV0_n, __A04_1__DV1, __A04_1__DV1_n, GND, __A04_1__DV376_n, __A04_1__DV376, NET_196, TL15, __A04_1__BR1, NET_215, VCC, SIM_RST);
    U74HC02 U4018(__A04_1__DV0, __A04_1__DIV_n, ST0_n, __A04_1__DV1, __A04_1__DIV_n, ST1_n, GND, __A04_1__DIV_n, ST4_n, __A04_1__DV4, __A04_1__DIV_n, __A04_1__ST376_n, __A04_1__DV376, VCC, SIM_RST);
    U74HC02 U4019(NET_182, SUMA16_n, SUMB16_n, NET_197, PHS4, PHS3_n, GND, UNF_n, TOV_n, NET_186, L15_n, NET_196, NET_191, VCC, SIM_RST);
    U74HC27 #(0, 0, 1) U4020(PHS4_n, WL16_n, NET_191, NET_187, NET_214, NET_194, GND, NET_193, NET_215, NET_190, NET_189, NET_187, TSGN_n, VCC, SIM_RST);
    U74HC02 U4021(NET_190, TSGN_n, PHS3_n, NET_189, NET_196, PHS3_n, GND, TOV_n, PHS2_n, NET_195, __A04_1__SGUM, NET_186, NET_185, VCC, SIM_RST);
    U74HC4002 U4022(NET_192, NET_182, PHS3_n, TSGU_n, PHS4, NET_183, GND, NET_184, WL16_n, WL15_n, WL14_n, WL13_n, NET_220, VCC, SIM_RST);
    U74LVC07 U4023(NET_185, NET_215, NET_194, NET_215, NET_193, NET_214, GND, NET_214, NET_188, NET_219, NET_220, NET_219, NET_218, VCC, SIM_RST);
    U74HC02 #(1, 0, 0, 0) U4024(NET_188, NET_195, NET_192, NET_200, TOV_n, OVF_n, GND, NET_211, PHS3_n, NET_206, TMZ_n, PHS4_n, NET_221, VCC, SIM_RST);
    U74HC04 U4025(NET_214, __A04_1__BR1_n, __A04_1__TSGN2, NET_211, NET_207, __A04_1__BR2, GND, BR2_n, NET_202, __A04_1__DV4_n, __A04_1__DV4, NET_324, NET_323, VCC, SIM_RST);
    U74HC27 U4026(GEQZRO_n, PHS4_n, WL16_n, PHS4_n, NET_211, NET_203, GND, NET_204, NET_203, NET_219, NET_202, NET_201, TPZG_n, VCC, SIM_RST);
    U74HC4002 U4027(NET_218, WL12_n, WL11_n, WL10_n, WL09_n, NET_225, GND, NET_224, WL08_n, WL07_n, WL06_n, WL05_n, NET_217, VCC, SIM_RST);
    U74HC4002 #(0, 1) U4028(NET_216, WL04_n, WL03_n, WL02_n, WL01_n, NET_227, GND, NET_226, NET_207, NET_206, NET_205, NET_195, NET_202, VCC, SIM_RST);
    wire U4029_12_NC;
    wire U4029_13_NC;
    U74LVC07 U4029(NET_217, NET_219, NET_216, NET_219, NET_221, NET_219, GND, NET_207, NET_199, NET_207, NET_204, U4029_12_NC, U4029_13_NC, VCC, SIM_RST);
    U74HC02 U4030(NET_205, TMZ_n, PHS3_n, NET_199, NET_201, NET_200, GND, SQ0_n, EXST0_n, NET_323, QC3_n, SQEXT_n, NET_277, VCC, SIM_RST);
    U74HC27 U4031(NET_324, SQR10, QC0_n, NET_324, SQR10_n, __A04_2__WRITE0, GND, __A04_2__RAND0, SQR10, NET_324, QC1_n, __A04_2__READ0, QC0_n, VCC, SIM_RST);
    U74HC04 U4032(__A04_2__READ0, __A04_2__READ0_n, __A04_2__WRITE0, __A04_2__WRITE0_n, __A04_2__WOR0, __A04_2__WOR0_n, GND, __A04_2__RXOR0_n, RXOR0, __A04_2__RUPT0_n, __A04_2__RUPT0, __A04_2__RUPT1_n, __A04_2__RUPT1, VCC, SIM_RST);
    U74HC27 U4033(QC1_n, SQR10_n, SQR10, NET_324, QC2_n, __A04_2__ROR0, GND, __A04_2__WOR0, QC2_n, NET_324, SQR10_n, __A04_2__WAND0, NET_324, VCC, SIM_RST);
    U74HC27 U4034(SQR10, NET_324, QC3_n, NET_324, SQR10_n, __A04_2__RUPT0, GND, NET_278, ST0_n, SQR12_n, SQ2_n, RXOR0, QC3_n, VCC, SIM_RST);
    U74HC04 U4035(NET_278, NET_276, __A04_2__INOUT, __A04_2__INOUT_n, NET_283, NET_308, GND, __A04_2__BR1B2_n, __A04_2__BR1B2, __A04_2__BR12B_n, __A04_2__BR12B, __A04_2__BR1B2B_n, BR1B2B, VCC, SIM_RST);
    U74HC02 U4036(__A04_2__PRINC, NET_277, NET_276, __A04_2__RRPA, T03_n, __A04_2__RUPT1_n, GND, T03_n, __A04_2__RXOR0_n, __A04_2__3XP7, NET_271, T03_n, NET_274, VCC, SIM_RST);
    U74HC27 U4037(EXST0_n, SQ0_n, __A04_2__INOUT, __A04_1__DV4, __A04_2__PRINC, __A04_2__8PP4, GND, NET_320, NET_274, NET_272, NET_279, __A04_2__INOUT, __A04_2__RUPT0_n, VCC, SIM_RST);
    U74HC02 U4038(NET_271, __A04_2__ROR0, __A04_2__WOR0, NET_273, T03_n, NET_275, GND, __A04_2__RAND0, __A04_2__WAND0, NET_275, __A04_1__DV4_n, T05_n, __A04_2__5XP28, VCC, SIM_RST);
    U74LVC07 U4039(NET_320, __A04_2__RB_n, NET_318, __A04_2__RC_n, NET_319, __A04_2__5XP11, GND, __A04_2__5XP11, NET_321, __A04_2__RA_n, NET_322, __A04_2__WG_n, NET_330, VCC, SIM_RST);
    U74HC27 U4040(NET_273, NET_287, T05_n, __A04_2__INOUT_n, __A04_2__READ0, NET_319, GND, __A04_2__WCH_n, NET_285, n7XP14, NET_286, NET_318, NET_281, VCC, SIM_RST);
    U74HC02 U4041(NET_321, __A04_2__WRITE0, RXOR0, NET_272, __A04_2__READ0_n, T05_n, GND, __A04_2__WRITE0_n, T05_n, NET_285, T05_n, __A04_2__WOR0_n, NET_286, VCC, SIM_RST);
    U74HC02 U4042(NET_287, T05_n, __A04_2__RXOR0_n, NET_280, T02_n, __A04_2__WRITE0_n, GND, T02_n, __A04_2__INOUT_n, __A04_2__2XP3, T09_n, __A04_2__RUPT0_n, __A04_2__9XP1, VCC, SIM_RST);
    U74HC27 U4043(NET_285, NET_287, __A04_2__RUPT1, IC13, IC12, NET_282, GND, NET_330, __A04_2__9XP1, NET_281, NET_279, NET_322, __A04_2__2XP3, VCC, SIM_RST);
    U74HC02 U4044(NET_281, T09_n, __A04_2__RXOR0_n, NET_279, T09_n, NET_282, GND, NET_287, NET_280, NET_329, T01_n, __A04_2__RUPT1_n, __A04_2__RB2, VCC, SIM_RST);
    U74LVC07 U4045(NET_329, __A04_2__WG_n, NET_328, NET_283, NET_327, NET_283, GND, __A04_2__RA_n, NET_305, __A04_2__WG_n, NET_314, TMZ_n, NET_317, VCC, SIM_RST);
    U74HC27 U4046(__A04_2__RUPT0, __A04_2__RUPT1, __A04_2__INOUT, MP1, MP3A, NET_328, GND, NET_327, __A04_1__DV0, IC15, __A04_1__DV1376, NET_284, RSM3, VCC, SIM_RST);
    U74HC02 U4047(__A04_2__R15, NET_284, T01_n, __A04_2__1XP10, T01_n, __A04_2__DV0_n, GND, MP0_n, T03_n, NET_301, __A04_2__INOUT_n, T03_n, NET_312, VCC, SIM_RST);
    U74HC27 U4048(T02_n, __A04_2__DV0_n, __A04_2__BRDIF_n, TS0_n, T04_n, NET_291, GND, NET_288, T04_n, __A04_1__BR1, MP0_n, __A04_2__2XP5, __A04_1__BR1, VCC, SIM_RST);
    U74HC02 U4049(__A04_2__3XP2, T03_n, TS0_n, __A04_2__BR1B2, __A04_1__BR1, BR2_n, GND, __A04_1__BR1_n, __A04_1__BR2, __A04_2__BR12B, __A04_2__BR1B2, __A04_2__BR12B, __A04_2__BRDIF_n, VCC, SIM_RST);
    U74HC02 U4050(BR1B2B, __A04_1__BR2, __A04_1__BR1, __A04_2__4XP5, TS0_n, T04_n, GND, T04_n, __A04_2__INOUT_n, __A04_2__4XP11, T04_n, MP3_n, NET_313, VCC, SIM_RST);
    U74HC27 U4051(MP0_n, __A04_1__BR1_n, __A04_1__DV1_n, T04_n, BR2_n, NET_302, GND, NET_296, TS0_n, T05_n, __A04_2__BR1B2_n, NET_269, T04_n, VCC, SIM_RST);
    U74HC27 U4052(T05_n, TS0_n, T07_n, __A04_1__BR1_n, MP3_n, __A04_2__7XP19, GND, __A04_2__8XP6, T08_n, __A04_1__DV1_n, __A04_1__BR2, NET_297, __A04_2__BR12B_n, VCC, SIM_RST);
    U74HC02 U4053(__A04_2__B15X, T05_n, __A04_1__DV1_n, n5XP4, T05_n, RSM3_n, GND, T06_n, __A04_1__DV1_n, __A04_2__6XP5, T06_n, MP3_n, TL15, VCC, SIM_RST);
    U74HC02 U4054(__A04_1__TSGN2, T07_n, MP0_n, NET_306, T07_n, __A04_1__DV1_n, GND, T08_n, __A04_1__DV1_n, __A04_2__8XP5, T09_n, MP3_n, NET_304, VCC, SIM_RST);
    U74HC27 U4055(T09_n, __A04_1__BR1, T09_n, MP0_n, __A04_1__BR1_n, NET_290, GND, NET_293, MP0_n, T09_n, __A04_2__BRDIF_n, NET_310, MP0_n, VCC, SIM_RST);
    U74HC02 U4056(KRPT, T09_n, __A04_2__RUPT1_n, __A04_2__MP0T10, T10_n, MP0_n, GND, NET_308, T02_n, NET_315, STORE1_n, T09_n, NET_316, VCC, SIM_RST);
    U74HC27 U4057(MP3_n, MP0_n, __A04_2__1XP10, __A04_2__8XP5, NET_304, NET_305, GND, __A04_2__RSC_n, NET_315, NET_313, NET_306, NET_307, T11_n, VCC, SIM_RST);
    wire U4058_8_NC;
    wire U4058_9_NC;
    wire U4058_10_NC;
    wire U4058_11_NC;
    wire U4058_12_NC;
    wire U4058_13_NC;
    U74HC04 U4058(__A04_2__RSC_n, __A04_2__MRSC, NET_307, NET_299, TRSM, NET_210, GND, U4058_8_NC, U4058_9_NC, U4058_10_NC, U4058_11_NC, U4058_12_NC, U4058_13_NC, VCC, SIM_RST);
    U74HC27 U4059(NET_315, NET_316, NET_312, __A04_2__B15X, __A04_2__7XP19, NET_309, GND, NET_311, __A04_2__8XP5, NET_310, NET_290, NET_314, NET_313, VCC, SIM_RST);
    U74HC02 U4060(NET_317, __A04_2__2XP5, __A04_2__1XP10, NET_292, NET_291, NET_293, GND, __A04_2__1XP10, __A04_2__MP0T10, NET_300, NET_296, NET_307, NET_298, VCC, SIM_RST);
    U74LVC07 U4061(NET_309, __A04_2__WY_n, NET_311, __A04_2__WY_n, NET_294, __A04_2__WL_n, GND, __A04_2__RC_n, NET_295, __A04_2__RB_n, NET_289, __A04_2__CI_n, NET_292, VCC, SIM_RST);
    U74HC27 U4062(NET_288, NET_269, NET_269, __A04_2__2XP5, NET_290, NET_295, GND, NET_289, NET_288, __A04_2__7XP19, NET_310, NET_294, __A04_2__6XP5, VCC, SIM_RST);
    wire U4063_10_NC;
    wire U4063_11_NC;
    wire U4063_12_NC;
    wire U4063_13_NC;
    U74LVC07 U4063(NET_300, TSGN_n, NET_303, TSGN_n, NET_298, __A04_2__RB1_n, GND, __A04_2__L16_n, NET_299, U4063_10_NC, U4063_11_NC, U4063_12_NC, U4063_13_NC, VCC, SIM_RST);
    wire U4064_3_NC;
    wire U4064_4_NC;
    wire U4064_5_NC;
    wire U4064_6_NC;
    wire U4064_8_NC;
    wire U4064_9_NC;
    wire U4064_10_NC;
    wire U4064_11_NC;
    U74HC27 U4064(NET_302, NET_301, U4064_3_NC, U4064_4_NC, U4064_5_NC, U4064_6_NC, GND, U4064_8_NC, U4064_9_NC, U4064_10_NC, U4064_11_NC, NET_303, NET_306, VCC, SIM_RST);
    wire U4065_4_NC;
    wire U4065_5_NC;
    wire U4065_6_NC;
    wire U4065_8_NC;
    wire U4065_9_NC;
    wire U4065_10_NC;
    wire U4065_11_NC;
    wire U4065_12_NC;
    wire U4065_13_NC;
    U74HC02 U4065(__A04_2__R1C_n, NET_307, NET_297, U4065_4_NC, U4065_5_NC, U4065_6_NC, GND, U4065_8_NC, U4065_9_NC, U4065_10_NC, U4065_11_NC, U4065_12_NC, U4065_13_NC, VCC, SIM_RST);
endmodule