`include "components/agc_parts.v"

module timer(VCC, GND, SIM_RST, CLOCK, MSTRTP, MSTP, PHS2, PHS2_n, PHS3_n, PHS4, PHS4_n, RT, RT_n, WT, WT_n, CT, CT_n, CLK, TT_n, P01, P01_n, P02, P02_n, P03, P03_n, P04, P04_n, P05, P05_n, SBY, ALGA, STRT1, STRT2, GOJ1, STOPA, GOJAM, GOJAM_n, STOP, STOP_n, MONWT, Q2A, MGOJAM, MSTPIT_n);
    input wire SIM_RST;
    wire __A02_1__cdiv_1__A;
    wire __A02_1__cdiv_2__C;
    wire __A02_1__cdiv_2__F;
    input wire GOJ1;
    wire __A02_1__oddset;
    output wire RT_n;
    output wire P02_n;
    output wire WT_n;
    wire NET_88;
    wire __A02_1__RINGA_n;
    wire NET_82;
    output wire MONWT;
    wire __A02_2__F01C;
    wire NET_85;
    output wire STOPA;
    wire NET_95;
    output wire GOJAM_n;
    wire __A02_1__cdiv_2__D;
    wire __A02_2__F01D;
    wire NET_76;
    output wire GOJAM;
    output wire P01;
    output wire PHS2_n;
    wire __A02_1__cdiv_2__FS;
    output wire P03;
    input wire VCC;
    wire __A02_1__ODDSET_n;
    input wire STRT2;
    wire __A02_2__FS01_n;
    wire __A02_1__RINGB_n;
    output wire STOP;
    wire __A02_1__ovfstb_r5;
    wire NET_81;
    output wire P03_n;
    output wire CT;
    wire __A02_1__ovfstb_r6;
    output wire P05_n;
    wire __A02_2__F01A;
    wire __A02_1__ovfstb_r4;
    wire __A02_1__ovfstb_r1;
    wire NET_90;
    wire NET_77;
    wire NET_97;
    input wire CLOCK;
    wire NET_79;
    wire NET_91;
    wire NET_75;
    output wire P01_n;
    input wire STRT1;
    output wire PHS4_n;
    wire NET_89;
    input wire SBY;
    output wire Q2A;
    wire __A02_2__FS01;
    wire __A02_1__cdiv_1__B;
    output wire P04;
    wire NET_94;
    output wire CT_n;
    wire __A02_1__cdiv_2__A;
    wire NET_83;
    input wire GND;
    wire __A02_1__OVFSTB_n;
    output wire MSTPIT_n;
    output wire CLK;
    output wire TT_n;
    wire __A02_1__cdiv_2__B;
    wire __A02_1__cdiv_2__FS_n;
    output wire P05;
    wire __A02_1__ovfstb_r2;
    wire NET_93;
    output wire PHS3_n;
    output wire P04_n;
    wire __A02_1__cdiv_1__FS;
    output wire STOP_n;
    output wire MGOJAM;
    wire __A02_1__evnset;
    wire NET_80;
    wire NET_96;
    output wire PHS2;
    input wire ALGA;
    output wire RT;
    input wire MSTRTP;
    wire NET_87;
    wire NET_84;
    output wire WT;
    wire __A02_1__cdiv_1__D;
    input wire MSTP;
    wire __A02_1__ovfstb_r3;
    wire __A02_2__F01B;
    output wire P02;
    wire NET_86;
    wire NET_61;
    output wire PHS4;
    wire __A02_1__cdiv_1__FS_n;
    wire __A02_1__EVNSET_n;
    wire NET_78;
    wire NET_92;

    U74HC04 U3(__A02_1__cdiv_1__D, __A02_1__cdiv_2__F, PHS2, PHS2_n, PHS4, PHS4_n, GND, NET_61, __A02_1__cdiv_1__B, CT, NET_61, CT_n, CT, VCC, SIM_RST);
    wire U7_8_NC;
    wire U7_9_NC;
    wire U7_10_NC;
    wire U7_11_NC;
    U74HC27 #(0, 1, 0) U7(__A02_1__cdiv_2__D, __A02_1__cdiv_2__F, __A02_1__cdiv_2__B, __A02_1__cdiv_2__F, __A02_1__cdiv_2__C, __A02_1__cdiv_2__A, GND, U7_8_NC, U7_9_NC, U7_10_NC, U7_11_NC, __A02_1__cdiv_2__B, __A02_1__cdiv_2__A, VCC, SIM_RST);
    wire U2_8_NC;
    wire U2_9_NC;
    wire U2_10_NC;
    wire U2_11_NC;
    U74HC27 #(0, 1, 0) U2(__A02_1__cdiv_1__D, CLOCK, __A02_1__cdiv_1__B, CLOCK, PHS2, __A02_1__cdiv_1__A, GND, U2_8_NC, U2_9_NC, U2_10_NC, U2_11_NC, __A02_1__cdiv_1__B, __A02_1__cdiv_1__A, VCC, SIM_RST);
    wire U4_8_NC;
    wire U4_9_NC;
    wire U4_10_NC;
    wire U4_11_NC;
    wire U4_12_NC;
    wire U4_13_NC;
    U74HC02 U4(PHS4, __A02_1__cdiv_2__F, __A02_1__cdiv_1__A, __A02_1__oddset, STOP, __A02_1__RINGA_n, GND, U4_8_NC, U4_9_NC, U4_10_NC, U4_11_NC, U4_12_NC, U4_13_NC, VCC, SIM_RST);
    U74HC27 U11(__A02_1__RINGB_n, P05_n, P04, P05, __A02_1__RINGA_n, NET_82, GND, NET_90, GND, NET_95, __A02_1__EVNSET_n, NET_83, P04_n, VCC, SIM_RST);
    U74HC04 U5(__A02_1__cdiv_1__FS_n, WT, WT, WT_n, WT, TT_n, GND, __A02_1__ovfstb_r5, __A02_1__ovfstb_r4, __A02_1__ovfstb_r6, __A02_1__ovfstb_r5, __A02_1__OVFSTB_n, __A02_1__ovfstb_r2, VCC, SIM_RST);
    U74HC02 U23(NET_91, NET_90, STOPA, STOPA, NET_91, NET_89, GND, NET_97, NET_94, NET_88, NET_88, NET_92, NET_94, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U15(P04, NET_76, P04_n, P04_n, P04, NET_77, GND, __A02_1__RINGB_n, P04, NET_81, P04_n, __A02_1__RINGA_n, NET_80, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U12(P01, NET_83, P01_n, P01_n, P01, NET_82, GND, __A02_1__RINGA_n, P01, NET_84, P01_n, __A02_1__RINGB_n, NET_78, VCC, SIM_RST);
    pullup R1(NET_95);
    U74HC04 U8(__A02_1__cdiv_2__D, __A02_1__RINGA_n, __A02_1__oddset, __A02_1__ODDSET_n, __A02_1__cdiv_2__C, __A02_1__RINGB_n, GND, __A02_1__evnset, __A02_1__RINGB_n, __A02_1__EVNSET_n, __A02_1__evnset, RT, __A02_1__cdiv_1__A, VCC, SIM_RST);
    U74HC02 #(0, 1, 1, 0) U16(P05, NET_81, P05_n, P05_n, P05, NET_80, GND, NET_95, GOJ1, NET_87, __A02_1__EVNSET_n, NET_96, NET_89, VCC, SIM_RST);
    U74HC27 U19(SBY, ALGA, STRT1, STRT2, NET_87, NET_85, GND, NET_97, GND, NET_93, __A02_1__EVNSET_n, NET_86, MSTRTP, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U17(__A02_2__F01D, __A02_2__FS01_n, __A02_2__F01B, __A02_2__FS01_n, __A02_2__F01B, __A02_2__FS01, GND, __A02_2__FS01_n, __A02_2__F01A, __A02_2__FS01, __A02_2__F01A, __A02_2__FS01, __A02_2__F01C, VCC, SIM_RST);
    wire U22_11_NC;
    wire U22_12_NC;
    wire U22_13_NC;
    U74HC02 U22(NET_92, __A02_1__EVNSET_n, MSTP, GOJAM_n, STRT2, STOPA, GND, STOPA, NET_94, STOP_n, U22_11_NC, U22_12_NC, U22_13_NC, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U6(__A02_1__cdiv_2__D, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__FS, GND, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__A, __A02_1__cdiv_2__FS, __A02_1__cdiv_2__A, __A02_1__cdiv_2__FS, __A02_1__cdiv_2__C, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U13(P02, NET_84, P02_n, P02_n, P02, NET_78, GND, __A02_1__RINGB_n, P02, NET_79, P02_n, __A02_1__RINGA_n, NET_75, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U1(__A02_1__cdiv_1__D, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__B, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__B, __A02_1__cdiv_1__FS, GND, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__A, __A02_1__cdiv_1__FS, __A02_1__cdiv_1__A, __A02_1__cdiv_1__FS, PHS2, VCC, SIM_RST);
    U74HC02 U9(__A02_1__ovfstb_r1, CT_n, __A02_1__ovfstb_r2, __A02_1__ovfstb_r2, __A02_1__ovfstb_r6, __A02_1__ovfstb_r1, GND, __A02_1__ovfstb_r4, __A02_1__ovfstb_r2, __A02_1__ovfstb_r3, __A02_1__ovfstb_r3, __A02_1__ovfstb_r1, __A02_1__ovfstb_r4, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U14(P03, NET_79, P03_n, P03_n, P03, NET_75, GND, __A02_1__RINGA_n, P03, NET_76, P03_n, __A02_1__RINGB_n, NET_77, VCC, SIM_RST);
    wire U18_8_NC;
    wire U18_9_NC;
    wire U18_10_NC;
    wire U18_11_NC;
    U74HC27 #(0, 1, 0) U18(__A02_2__F01D, P01_n, __A02_2__F01B, P01_n, __A02_2__F01C, __A02_2__F01A, GND, U18_8_NC, U18_9_NC, U18_10_NC, U18_11_NC, __A02_2__F01B, __A02_2__F01A, VCC, SIM_RST);
    U74HC04 U21(NET_95, NET_96, MSTP, NET_93, GOJAM_n, GOJAM, GND, MGOJAM, GOJAM, STOP, STOP_n, MSTPIT_n, STOP, VCC, SIM_RST);
    wire U10_12_NC;
    wire U10_13_NC;
    U74HC04 U10(CT, PHS3_n, WT_n, CLK, WT_n, MONWT, GND, Q2A, WT_n, RT_n, RT, U10_12_NC, U10_13_NC, VCC, SIM_RST);
    wire U20_5_NC;
    wire U20_6_NC;
    wire U20_8_NC;
    wire U20_9_NC;
    wire U20_10_NC;
    wire U20_11_NC;
    wire U20_12_NC;
    wire U20_13_NC;
    U74LVC07 U20(NET_86, NET_95, NET_85, NET_95, U20_5_NC, U20_6_NC, GND, U20_8_NC, U20_9_NC, U20_10_NC, U20_11_NC, U20_12_NC, U20_13_NC, VCC, SIM_RST);
endmodule