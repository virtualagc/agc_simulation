`timescale 1ns/1ps

module four_bit_2(VCC, GND, SIM_RST, A2XG_n, CAG, CBG, CGG, CLG1G, CLXC, CQG, CUG, CZG, L2GDG_n, RAG_n, RCG_n, RGG_n, RLG_n, RQG_n, RZG_n, WAG_n, WALSG_n, WBG_n, WLG_n, WQG_n, WZG_n, CI05_n, CO06, MONEX, XUY09_n, XUY10_n, CH05, CH06, CH07, CH08, G05ED, G06ED, G07ED, L04_n, G2LSG_n, G09_n, G10_n, G11_n, MDT05, MDT06, MDT07, MDT08, SA05, SA06, SA07, SA08, RBLG_n, RULOG_n, WL09_n, WL10_n, WG1G_n, WG3G_n, WG4G_n, WYDG_n, WYLOG_n, R1C, WL04_n, CI09_n, CO10, G05_n, G06_n, G07_n, L08_n, XUY05_n, XUY06_n, WL05_n, WL06_n, WL07_n, WL08_n);
    input wire SIM_RST;
    input wire A2XG_n;
    input wire CAG;
    input wire CBG;
    input wire CGG;
    input wire CH05;
    input wire CH06;
    input wire CH07;
    input wire CH08;
    input wire CI05_n;
    output wire CI09_n;
    input wire CLG1G;
    input wire CLXC;
    input wire CO06;
    inout wire CO10;
    input wire CQG;
    input wire CUG;
    input wire CZG;
    input wire G05ED;
    inout wire G05_n;
    input wire G06ED;
    inout wire G06_n;
    input wire G07ED;
    inout wire G07_n;
    input wire G09_n;
    input wire G10_n;
    input wire G11_n;
    input wire G2LSG_n;
    input wire GND;
    input wire L04_n;
    inout wire L08_n;
    input wire L2GDG_n;
    input wire MDT05;
    input wire MDT06;
    input wire MDT07;
    input wire MDT08;
    input wire MONEX;
    wire NET_125;
    wire NET_126;
    wire NET_127;
    wire NET_128;
    wire NET_129;
    wire NET_130;
    wire NET_131;
    wire NET_132;
    wire NET_133;
    wire NET_134;
    wire NET_135;
    wire NET_138;
    wire NET_139;
    wire NET_140;
    wire NET_141;
    wire NET_142;
    wire NET_143;
    wire NET_144;
    wire NET_148;
    wire NET_149;
    wire NET_150;
    wire NET_151;
    wire NET_152;
    wire NET_153;
    wire NET_154;
    wire NET_155;
    wire NET_156;
    wire NET_159;
    wire NET_160;
    wire NET_161;
    wire NET_162;
    wire NET_163;
    wire NET_164;
    wire NET_165;
    wire NET_166;
    wire NET_167;
    wire NET_168;
    wire NET_169;
    wire NET_170;
    wire NET_171;
    wire NET_172;
    wire NET_173;
    wire NET_174;
    wire NET_175;
    wire NET_176;
    wire NET_177;
    wire NET_178;
    wire NET_179;
    wire NET_180;
    wire NET_181;
    wire NET_182;
    wire NET_183;
    wire NET_184;
    wire NET_185;
    wire NET_190;
    wire NET_191;
    wire NET_192;
    wire NET_193;
    wire NET_194;
    wire NET_195;
    wire NET_196;
    wire NET_197;
    wire NET_198;
    wire NET_199;
    wire NET_200;
    wire NET_201;
    wire NET_202;
    wire NET_203;
    wire NET_204;
    wire NET_205;
    wire NET_206;
    wire NET_207;
    wire NET_208;
    wire NET_209;
    wire NET_210;
    wire NET_211;
    wire NET_212;
    wire NET_213;
    wire NET_214;
    wire NET_215;
    wire NET_216;
    wire NET_217;
    wire NET_218;
    wire NET_219;
    wire NET_220;
    wire NET_221;
    wire NET_222;
    wire NET_223;
    wire NET_224;
    wire NET_225;
    wire NET_226;
    wire NET_229;
    wire NET_230;
    wire NET_231;
    wire NET_232;
    wire NET_233;
    wire NET_234;
    wire NET_235;
    wire NET_239;
    wire NET_240;
    wire NET_241;
    wire NET_242;
    wire NET_243;
    wire NET_244;
    wire NET_245;
    wire NET_246;
    wire NET_247;
    wire NET_250;
    wire NET_251;
    wire NET_252;
    wire NET_253;
    wire NET_254;
    wire NET_255;
    wire NET_256;
    wire NET_257;
    wire NET_258;
    wire NET_259;
    wire NET_260;
    wire NET_261;
    wire NET_262;
    wire NET_263;
    wire NET_264;
    wire NET_265;
    wire NET_266;
    wire NET_267;
    wire NET_268;
    wire NET_269;
    wire NET_270;
    wire NET_271;
    wire NET_272;
    wire NET_273;
    wire NET_274;
    wire NET_275;
    wire NET_276;
    wire NET_281;
    wire NET_282;
    wire NET_283;
    wire NET_284;
    wire NET_285;
    wire NET_286;
    wire NET_287;
    wire NET_288;
    wire NET_289;
    wire NET_290;
    wire NET_291;
    wire NET_292;
    wire NET_293;
    wire NET_294;
    wire NET_295;
    wire NET_296;
    wire NET_297;
    wire NET_298;
    wire NET_299;
    wire NET_300;
    wire NET_301;
    wire NET_302;
    wire NET_303;
    wire NET_304;
    wire NET_305;
    wire NET_306;
    input wire R1C;
    input wire RAG_n;
    input wire RBLG_n;
    input wire RCG_n;
    input wire RGG_n;
    input wire RLG_n;
    input wire RQG_n;
    input wire RULOG_n;
    input wire RZG_n;
    input wire SA05;
    input wire SA06;
    input wire SA07;
    input wire SA08;
    input wire VCC;
    input wire WAG_n;
    input wire WALSG_n;
    input wire WBG_n;
    input wire WG1G_n;
    input wire WG3G_n;
    input wire WG4G_n;
    input wire WL04_n;
    output wire WL05_n;
    output wire WL06_n;
    output wire WL07_n;
    output wire WL08_n;
    input wire WL09_n;
    input wire WL10_n;
    input wire WLG_n;
    input wire WQG_n;
    input wire WYDG_n;
    input wire WYLOG_n;
    input wire WZG_n;
    output wire XUY05_n;
    output wire XUY06_n;
    input wire XUY09_n;
    input wire XUY10_n;
    wire __A09_1__X1;
    wire __A09_1__X1_n;
    wire __A09_1__X2;
    wire __A09_1__X2_n;
    wire __A09_1__Y1;
    wire __A09_1__Y1_n;
    wire __A09_1__Y2;
    wire __A09_1__Y2_n;
    wire __A09_1___A1_n;
    wire __A09_1___A2_n;
    wire __A09_1___B1_n;
    wire __A09_1___B2_n;
    wire __A09_1___CI_INTERNAL;
    wire __A09_1___G1;
    wire __A09_1___G2;
    wire __A09_1___GEM1;
    wire __A09_1___GEM2;
    wire __A09_1___L1_n;
    wire __A09_1___L2_n;
    wire __A09_1___MWL1;
    wire __A09_1___MWL2;
    wire __A09_1___Q1_n;
    wire __A09_1___Q2_n;
    wire __A09_1___RL1_n;
    wire __A09_1___RL2_n;
    wire __A09_1___SUMA1;
    wire __A09_1___SUMA2;
    wire __A09_1___SUMB1;
    wire __A09_1___SUMB2;
    wire __A09_1___WL1;
    wire __A09_1___WL2;
    wire __A09_1___Z1_n;
    wire __A09_1___Z2_n;
    wire __A09_2__X1;
    wire __A09_2__X1_n;
    wire __A09_2__X2;
    wire __A09_2__X2_n;
    wire __A09_2__Y1;
    wire __A09_2__Y1_n;
    wire __A09_2__Y2;
    wire __A09_2__Y2_n;
    wire __A09_2___A1_n;
    wire __A09_2___A2_n;
    wire __A09_2___B1_n;
    wire __A09_2___B2_n;
    wire __A09_2___CI_IN;
    wire __A09_2___CI_INTERNAL;
    wire __A09_2___CO_IN;
    wire __A09_2___G1;
    wire __A09_2___G2;
    wire __A09_2___G2_n;
    wire __A09_2___GEM1;
    wire __A09_2___GEM2;
    wire __A09_2___L1_n;
    wire __A09_2___MWL1;
    wire __A09_2___MWL2;
    wire __A09_2___Q1_n;
    wire __A09_2___Q2_n;
    wire __A09_2___RL1_n;
    wire __A09_2___RL2_n;
    wire __A09_2___SUMA1;
    wire __A09_2___SUMA2;
    wire __A09_2___SUMB1;
    wire __A09_2___SUMB2;
    wire __A09_2___WL1;
    wire __A09_2___WL2;
    wire __A09_2___XUY1;
    wire __A09_2___XUY2;
    wire __A09_2___Z1_n;
    wire __A09_2___Z2_n;

    pullup R9001(__A09_2___CO_IN);
    pullup R9002(__A09_1___RL1_n);
    pullup R9003(__A09_1___L1_n);
    pullup R9005(__A09_1___Z1_n);
    pullup R9006(G05_n);
    pullup R9007(__A09_1___RL2_n);
    pullup R9008(__A09_1___L2_n);
    pullup R9009(__A09_1___Z2_n);
    pullup R9010(G06_n);
    pullup R9011(CO10);
    pullup R9012(__A09_2___RL1_n);
    pullup R9013(__A09_2___L1_n);
    pullup R9015(__A09_2___Z1_n);
    pullup R9016(G07_n);
    pullup R9017(__A09_2___RL2_n);
    pullup R9018(L08_n);
    pullup R9019(__A09_2___Z2_n);
    pullup R9020(__A09_2___G2_n);
    U74HC02 U9001(NET_190, A2XG_n, __A09_1___A1_n, NET_185, WYLOG_n, WL05_n, GND, WL04_n, WYDG_n, NET_184, __A09_1__Y1_n, CUG, __A09_1__Y1, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U9002(MONEX, NET_190, __A09_1__X1_n, CLXC, CUG, __A09_1__X1, GND, __A09_1__Y1_n, NET_185, NET_184, __A09_1__Y1, __A09_1__X1_n, __A09_1__X1, VCC, SIM_RST);
    U74HC02 U9003(NET_193, __A09_1__X1_n, __A09_1__Y1_n, XUY05_n, __A09_1__X1, __A09_1__Y1, GND, NET_193, XUY05_n, NET_192, NET_193, __A09_1___SUMA1, __A09_1___CI_INTERNAL, VCC, SIM_RST);
    U74HC27 U9004(NET_193, XUY05_n, __A09_1___SUMA1, __A09_1___SUMB1, RULOG_n, NET_175, GND, NET_177, __A09_2___XUY1, XUY05_n, CI05_n, __A09_1___SUMA1, CI05_n, VCC, SIM_RST);
    U74HC04 U9005(CI05_n, NET_191, G05_n, __A09_1___GEM1, __A09_1___RL1_n, __A09_1___WL1, GND, WL05_n, __A09_1___WL1, __A09_1___MWL1, __A09_1___RL1_n, NET_138, __A09_1___CI_INTERNAL, VCC, SIM_RST);
    U74HC02 U9006(__A09_1___SUMB1, NET_192, NET_191, NET_176, WAG_n, WL05_n, GND, WL07_n, WALSG_n, NET_173, __A09_1___A1_n, CAG, NET_172, VCC, SIM_RST);
    U74LVC07 U9007(NET_177, __A09_2___CO_IN, NET_174, __A09_1___RL1_n, NET_183, __A09_1___L1_n, GND, __A09_1___Z1_n, NET_207, __A09_1___RL1_n, NET_208, __A09_1___RL1_n, NET_214, VCC, SIM_RST);
    U74HC02 U9008(NET_171, RAG_n, __A09_1___A1_n, NET_180, WLG_n, WL05_n, GND, __A09_2___G2_n, G2LSG_n, NET_182, __A09_1___L1_n, CLG1G, NET_181, VCC, SIM_RST);
    wire U9009_1_NC;
    wire U9009_2_NC;
    wire U9009_3_NC;
    U74HC02 #(0, 0, 1, 0) U9009(U9009_1_NC, U9009_2_NC, U9009_3_NC, NET_178, WQG_n, WL05_n, GND, NET_178, NET_179, __A09_1___Q1_n, __A09_1___Q1_n, CQG, NET_179, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U9010(NET_202, RQG_n, __A09_1___Q1_n, NET_210, WZG_n, WL05_n, GND, NET_210, NET_206, NET_207, __A09_1___Z1_n, CZG, NET_206, VCC, SIM_RST);
    U74HC27 U9011(NET_212, NET_202, MDT05, R1C, GND, NET_214, GND, NET_211, NET_198, NET_197, NET_203, NET_208, NET_209, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U9012(NET_209, RZG_n, __A09_1___Z1_n, NET_215, WBG_n, WL05_n, GND, NET_215, NET_213, __A09_1___B1_n, __A09_1___B1_n, CBG, NET_213, VCC, SIM_RST);
    U74LVC07 U9013(NET_140, __A09_2___CO_IN, NET_211, __A09_1___RL1_n, NET_194, G05_n, GND, G05_n, NET_195, __A09_1___RL2_n, NET_127, __A09_1___L2_n, NET_166, VCC, SIM_RST);
    U74HC02 U9014(NET_198, RBLG_n, __A09_1___B1_n, NET_197, NET_213, RCG_n, GND, WL04_n, WG3G_n, NET_201, WL06_n, WG4G_n, NET_200, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U9015(NET_176, NET_173, NET_175, NET_171, CH05, NET_174, GND, NET_183, NET_180, NET_182, NET_181, __A09_1___A1_n, NET_172, VCC, SIM_RST);
    U74HC02 U9016(NET_199, L2GDG_n, L04_n, NET_196, WG1G_n, WL05_n, GND, G05_n, CGG, __A09_1___G1, RGG_n, G05_n, NET_203, VCC, SIM_RST);
    wire U9017_3_NC;
    wire U9017_4_NC;
    wire U9017_5_NC;
    wire U9017_6_NC;
    U74HC27 #(1, 0, 0) U9017(NET_199, NET_196, U9017_3_NC, U9017_4_NC, U9017_5_NC, U9017_6_NC, GND, NET_212, RLG_n, __A09_1___L1_n, GND, NET_195, __A09_1___G1, VCC, SIM_RST);
    U74HC4002 U9018(NET_194, G05ED, SA05, NET_201, NET_200, NET_205, GND, NET_204, G06ED, SA06, NET_151, NET_150, NET_153, VCC, SIM_RST);
    U74HC02 U9019(NET_129, A2XG_n, __A09_1___A2_n, NET_143, WYLOG_n, WL06_n, GND, WL05_n, WYDG_n, NET_144, __A09_1__Y2_n, CUG, __A09_1__Y2, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U9020(MONEX, NET_129, __A09_1__X2_n, CLXC, CUG, __A09_1__X2, GND, __A09_1__Y2_n, NET_143, NET_144, __A09_1__Y2, __A09_1__X2_n, __A09_1__X2, VCC, SIM_RST);
    U74HC02 U9021(NET_141, __A09_1__X2_n, __A09_1__Y2_n, XUY06_n, __A09_1__X2, __A09_1__Y2, GND, __A09_2___XUY2, XUY06_n, NET_140, NET_141, XUY06_n, NET_139, VCC, SIM_RST);
    U74HC27 U9022(NET_141, XUY06_n, NET_141, __A09_1___SUMA2, CO06, __A09_2___CI_IN, GND, NET_142, __A09_1___SUMA2, __A09_1___SUMB2, RULOG_n, __A09_1___SUMA2, __A09_1___CI_INTERNAL, VCC, SIM_RST);
    U74HC02 U9023(__A09_1___SUMB2, NET_139, NET_138, NET_128, WAG_n, WL06_n, GND, WL08_n, WALSG_n, NET_130, __A09_1___A2_n, CAG, NET_126, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U9024(NET_128, NET_130, NET_142, NET_125, CH06, NET_127, GND, NET_166, NET_169, NET_170, NET_162, __A09_1___A2_n, NET_126, VCC, SIM_RST);
    U74HC02 U9025(NET_125, RAG_n, __A09_1___A2_n, NET_169, WLG_n, WL06_n, GND, G09_n, G2LSG_n, NET_170, __A09_1___L2_n, CLG1G, NET_162, VCC, SIM_RST);
    U74HC27 U9026(RLG_n, __A09_1___L2_n, NET_164, NET_163, NET_131, NET_132, GND, NET_135, MDT06, R1C, GND, NET_164, GND, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U9027(NET_160, WQG_n, WL06_n, __A09_1___Q2_n, NET_160, NET_161, GND, __A09_1___Q2_n, CQG, NET_161, RQG_n, __A09_1___Q2_n, NET_163, VCC, SIM_RST);
    U74LVC07 U9028(NET_132, __A09_1___RL2_n, NET_133, __A09_1___Z2_n, NET_135, __A09_1___RL2_n, GND, __A09_1___RL2_n, NET_156, G06_n, NET_153, G06_n, NET_152, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U9029(NET_165, WZG_n, WL06_n, NET_133, NET_165, NET_134, GND, __A09_1___Z2_n, CZG, NET_134, RZG_n, __A09_1___Z2_n, NET_131, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U9030(NET_167, WBG_n, WL06_n, __A09_1___B2_n, NET_167, NET_168, GND, __A09_1___B2_n, CBG, NET_168, RBLG_n, __A09_1___B2_n, NET_155, VCC, SIM_RST);
    wire U9031_8_NC;
    wire U9031_9_NC;
    wire U9031_10_NC;
    wire U9031_11_NC;
    U74HC27 #(0, 1, 0) U9031(NET_155, NET_154, NET_149, NET_148, __A09_1___G2, NET_152, GND, U9031_8_NC, U9031_9_NC, U9031_10_NC, U9031_11_NC, NET_156, NET_159, VCC, SIM_RST);
    U74HC02 U9032(NET_154, NET_168, RCG_n, NET_151, WL05_n, WG3G_n, GND, WL07_n, WG4G_n, NET_150, L2GDG_n, __A09_1___L1_n, NET_149, VCC, SIM_RST);
    wire U9033_11_NC;
    wire U9033_12_NC;
    wire U9033_13_NC;
    U74HC02 U9033(NET_148, WG1G_n, WL06_n, __A09_1___G2, G06_n, CGG, GND, RGG_n, G06_n, NET_159, U9033_11_NC, U9033_12_NC, U9033_13_NC, VCC, SIM_RST);
    wire U9034_10_NC;
    wire U9034_11_NC;
    wire U9034_12_NC;
    wire U9034_13_NC;
    U74HC04 U9034(G06_n, __A09_1___GEM2, __A09_1___RL2_n, __A09_1___WL2, __A09_1___WL2, WL06_n, GND, __A09_1___MWL2, __A09_1___RL2_n, U9034_10_NC, U9034_11_NC, U9034_12_NC, U9034_13_NC, VCC, SIM_RST);
    U74HC02 U9035(NET_281, A2XG_n, __A09_2___A1_n, NET_276, WYLOG_n, WL07_n, GND, WL06_n, WYDG_n, NET_275, __A09_2__Y1_n, CUG, __A09_2__Y1, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U9036(MONEX, NET_281, __A09_2__X1_n, CLXC, CUG, __A09_2__X1, GND, __A09_2__Y1_n, NET_276, NET_275, __A09_2__Y1, __A09_2__X1_n, __A09_2__X1, VCC, SIM_RST);
    U74HC02 U9037(NET_284, __A09_2__X1_n, __A09_2__Y1_n, __A09_2___XUY1, __A09_2__X1, __A09_2__Y1, GND, NET_284, __A09_2___XUY1, NET_283, NET_284, __A09_2___SUMA1, __A09_2___CI_INTERNAL, VCC, SIM_RST);
    U74HC27 U9038(NET_284, __A09_2___XUY1, __A09_2___SUMA1, __A09_2___SUMB1, RULOG_n, NET_266, GND, NET_268, XUY09_n, __A09_2___XUY1, __A09_2___CI_IN, __A09_2___SUMA1, __A09_2___CI_IN, VCC, SIM_RST);
    U74HC04 U9039(__A09_2___CI_IN, NET_282, G07_n, __A09_2___GEM1, __A09_2___RL1_n, __A09_2___WL1, GND, WL07_n, __A09_2___WL1, __A09_2___MWL1, __A09_2___RL1_n, NET_229, __A09_2___CI_INTERNAL, VCC, SIM_RST);
    U74HC02 U9040(__A09_2___SUMB1, NET_283, NET_282, NET_267, WAG_n, WL07_n, GND, WL09_n, WALSG_n, NET_264, __A09_2___A1_n, CAG, NET_263, VCC, SIM_RST);
    U74LVC07 U9041(NET_268, CO10, NET_265, __A09_2___RL1_n, NET_274, __A09_2___L1_n, GND, __A09_2___Z1_n, NET_298, __A09_2___RL1_n, NET_299, __A09_2___RL1_n, NET_305, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U9042(NET_267, NET_264, NET_266, NET_262, CH07, NET_265, GND, NET_274, NET_271, NET_273, NET_272, __A09_2___A1_n, NET_263, VCC, SIM_RST);
    U74HC02 U9043(NET_262, RAG_n, __A09_2___A1_n, NET_271, WLG_n, WL07_n, GND, G10_n, G2LSG_n, NET_273, __A09_2___L1_n, CLG1G, NET_272, VCC, SIM_RST);
    wire U9044_1_NC;
    wire U9044_2_NC;
    wire U9044_3_NC;
    wire U9044_4_NC;
    wire U9044_5_NC;
    wire U9044_6_NC;
    wire U9044_12_NC;
    wire U9044_13_NC;
    U74HC27 U9044(U9044_1_NC, U9044_2_NC, U9044_3_NC, U9044_4_NC, U9044_5_NC, U9044_6_NC, GND, NET_302, RLG_n, __A09_2___L1_n, GND, U9044_12_NC, U9044_13_NC, VCC, SIM_RST);
    wire U9045_1_NC;
    wire U9045_2_NC;
    wire U9045_3_NC;
    U74HC02 #(0, 0, 1, 0) U9045(U9045_1_NC, U9045_2_NC, U9045_3_NC, NET_269, WQG_n, WL07_n, GND, NET_269, NET_270, __A09_2___Q1_n, __A09_2___Q1_n, CQG, NET_270, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U9046(NET_285, RQG_n, __A09_2___Q1_n, NET_301, WZG_n, WL07_n, GND, NET_301, NET_297, NET_298, __A09_2___Z1_n, CZG, NET_297, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U9047(NET_300, RZG_n, __A09_2___Z1_n, NET_306, WBG_n, WL07_n, GND, NET_306, NET_304, __A09_2___B1_n, __A09_2___B1_n, CBG, NET_304, VCC, SIM_RST);
    U74HC02 U9048(NET_290, RBLG_n, __A09_2___B1_n, NET_289, NET_304, RCG_n, GND, WL06_n, WG3G_n, NET_293, WL08_n, WG4G_n, NET_292, VCC, SIM_RST);
    U74HC27 U9049(NET_302, NET_285, MDT07, R1C, GND, NET_305, GND, NET_303, NET_290, NET_289, NET_294, NET_299, NET_300, VCC, SIM_RST);
    U74LVC07 U9050(NET_231, CO10, NET_303, __A09_2___RL1_n, NET_286, G07_n, GND, G07_n, NET_287, __A09_2___RL2_n, NET_218, L08_n, NET_257, VCC, SIM_RST);
    U74HC02 U9051(NET_291, L2GDG_n, __A09_1___L2_n, NET_288, WG1G_n, WL07_n, GND, G07_n, CGG, __A09_2___G1, RGG_n, G07_n, NET_294, VCC, SIM_RST);
    U74HC4002 U9052(NET_286, G07ED, SA07, NET_293, NET_292, NET_296, GND, NET_295, GND, SA08, NET_242, NET_241, NET_244, VCC, SIM_RST);
    wire U9053_3_NC;
    wire U9053_4_NC;
    wire U9053_5_NC;
    wire U9053_6_NC;
    wire U9053_8_NC;
    wire U9053_9_NC;
    wire U9053_10_NC;
    wire U9053_11_NC;
    U74HC27 #(1, 0, 0) U9053(NET_291, NET_288, U9053_3_NC, U9053_4_NC, U9053_5_NC, U9053_6_NC, GND, U9053_8_NC, U9053_9_NC, U9053_10_NC, U9053_11_NC, NET_287, __A09_2___G1, VCC, SIM_RST);
    U74HC02 U9054(NET_220, A2XG_n, __A09_2___A2_n, NET_234, WYLOG_n, WL08_n, GND, WL07_n, WYDG_n, NET_235, __A09_2__Y2_n, CUG, __A09_2__Y2, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U9055(MONEX, NET_220, __A09_2__X2_n, CLXC, CUG, __A09_2__X2, GND, __A09_2__Y2_n, NET_234, NET_235, __A09_2__Y2, __A09_2__X2_n, __A09_2__X2, VCC, SIM_RST);
    U74HC02 U9056(NET_232, __A09_2__X2_n, __A09_2__Y2_n, __A09_2___XUY2, __A09_2__X2, __A09_2__Y2, GND, XUY10_n, __A09_2___XUY2, NET_231, NET_232, __A09_2___XUY2, NET_230, VCC, SIM_RST);
    U74HC27 U9057(NET_232, __A09_2___XUY2, NET_232, __A09_2___SUMA2, __A09_2___CO_IN, CI09_n, GND, NET_233, __A09_2___SUMA2, __A09_2___SUMB2, RULOG_n, __A09_2___SUMA2, __A09_2___CI_INTERNAL, VCC, SIM_RST);
    U74HC02 U9058(__A09_2___SUMB2, NET_230, NET_229, NET_219, WAG_n, WL08_n, GND, WL10_n, WALSG_n, NET_221, __A09_2___A2_n, CAG, NET_217, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U9059(NET_219, NET_221, NET_233, NET_216, CH08, NET_218, GND, NET_257, NET_260, NET_261, NET_253, __A09_2___A2_n, NET_217, VCC, SIM_RST);
    U74HC02 U9060(NET_216, RAG_n, __A09_2___A2_n, NET_260, WLG_n, WL08_n, GND, G11_n, G2LSG_n, NET_261, L08_n, CLG1G, NET_253, VCC, SIM_RST);
    U74HC27 U9061(RLG_n, L08_n, NET_255, NET_254, NET_222, NET_223, GND, NET_226, MDT08, R1C, GND, NET_255, GND, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U9062(NET_251, WQG_n, WL08_n, __A09_2___Q2_n, NET_251, NET_252, GND, __A09_2___Q2_n, CQG, NET_252, RQG_n, __A09_2___Q2_n, NET_254, VCC, SIM_RST);
    U74LVC07 U9063(NET_223, __A09_2___RL2_n, NET_224, __A09_2___Z2_n, NET_226, __A09_2___RL2_n, GND, __A09_2___RL2_n, NET_247, __A09_2___G2_n, NET_244, __A09_2___G2_n, NET_243, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U9064(NET_256, WZG_n, WL08_n, NET_224, NET_256, NET_225, GND, __A09_2___Z2_n, CZG, NET_225, RZG_n, __A09_2___Z2_n, NET_222, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U9065(NET_258, WBG_n, WL08_n, __A09_2___B2_n, NET_258, NET_259, GND, __A09_2___B2_n, CBG, NET_259, RBLG_n, __A09_2___B2_n, NET_246, VCC, SIM_RST);
    wire U9066_8_NC;
    wire U9066_9_NC;
    wire U9066_10_NC;
    wire U9066_11_NC;
    U74HC27 #(0, 1, 0) U9066(NET_246, NET_245, NET_240, NET_239, __A09_2___G2, NET_243, GND, U9066_8_NC, U9066_9_NC, U9066_10_NC, U9066_11_NC, NET_247, NET_250, VCC, SIM_RST);
    U74HC02 U9067(NET_245, NET_259, RCG_n, NET_242, WL07_n, WG3G_n, GND, WL09_n, WG4G_n, NET_241, L2GDG_n, __A09_2___L1_n, NET_240, VCC, SIM_RST);
    wire U9068_11_NC;
    wire U9068_12_NC;
    wire U9068_13_NC;
    U74HC02 U9068(NET_239, WG1G_n, WL08_n, __A09_2___G2, __A09_2___G2_n, CGG, GND, RGG_n, __A09_2___G2_n, NET_250, U9068_11_NC, U9068_12_NC, U9068_13_NC, VCC, SIM_RST);
    wire U9069_10_NC;
    wire U9069_11_NC;
    wire U9069_12_NC;
    wire U9069_13_NC;
    U74HC04 U9069(__A09_2___G2_n, __A09_2___GEM2, __A09_2___RL2_n, __A09_2___WL2, __A09_2___WL2, WL08_n, GND, __A09_2___MWL2, __A09_2___RL2_n, U9069_10_NC, U9069_11_NC, U9069_12_NC, U9069_13_NC, VCC, SIM_RST);
endmodule