`timescale 1ns/1ps
`default_nettype none

module four_bit_4(SIM_RST, SIM_CLK, p4VSW, GND, A2XG_n, CAG, CBG, CGG, CLG1G, CLG2G, CLXC, CQG, CUG, CZG, L2GDG_n, RAG_n, RCG_n, RGG_n, RLG_n, RQG_n, RZG_n, WAG_n, WALSG_n, WBG_n, WLG_n, WQG_n, WZG_n, CI13_n, CO14, BXVX, MONEX, XUY01_n, XUY02_n, CH13, CH14, CH16, L12_n, L16_n, G2LSG_n, WL01_n, WL02_n, G01_n, MDT13, MDT14, MDT15, MDT16, SA13, SA14, SA16, RBHG_n, RULOG_n, RUG_n, G16SW_n, WG1G_n, WG2G_n, WG3G_n, WG4G_n, WG5G_n, WYDG_n, WYHIG_n, R1C, US2SG, WL12_n, WHOMPA, Z15_n, Z16_n, A15_n, A16_n, EAC_n, G13, G13_n, G14, G14_n, G15, G15_n, G16, L15_n, RL13_n, RL14_n, RL15_n, RL16_n, SUMA13_n, SUMB13_n, SUMA14_n, SUMB14_n, SUMA15_n, SUMB15_n, SUMA16_n, SUMB16_n, WL13, WL13_n, WL14, WL14_n, WL15, WL15_n, WL16, WL16_n, XUY13_n, XUY14_n, GEM13, GEM14, GEM16, MWL13, MWL14, MWL15, MWL16);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    output wire A15_n;
    output wire A16_n;
    input wire A2XG_n;
    input wire BXVX;
    input wire CAG;
    input wire CBG;
    input wire CGG;
    input wire CH13;
    input wire CH14;
    input wire CH16;
    input wire CI13_n;
    input wire CLG1G;
    input wire CLG2G;
    input wire CLXC;
    input wire CO14;
    input wire CQG;
    input wire CUG;
    input wire CZG;
    output wire EAC_n;
    input wire G01_n;
    output wire G13;
    inout wire G13_n; //FPGA#wand
    output wire G14;
    inout wire G14_n; //FPGA#wand
    output wire G15;
    inout wire G15_n; //FPGA#wand
    output wire G16;
    input wire G16SW_n;
    input wire G2LSG_n;
    output wire GEM13;
    output wire GEM14;
    output wire GEM16;
    input wire L12_n;
    inout wire L15_n; //FPGA#wand
    inout wire L16_n; //FPGA#wand
    input wire L2GDG_n;
    input wire MDT13;
    input wire MDT14;
    input wire MDT15;
    input wire MDT16;
    input wire MONEX;
    output wire MWL13;
    output wire MWL14;
    output wire MWL15;
    output wire MWL16;
    input wire R1C;
    input wire RAG_n;
    input wire RBHG_n;
    input wire RCG_n;
    input wire RGG_n;
    inout wire RL13_n; //FPGA#wand
    inout wire RL14_n; //FPGA#wand
    inout wire RL15_n; //FPGA#wand
    inout wire RL16_n; //FPGA#wand
    input wire RLG_n;
    input wire RQG_n;
    input wire RUG_n;
    input wire RULOG_n;
    input wire RZG_n;
    input wire SA13;
    input wire SA14;
    input wire SA16;
    output wire SUMA13_n;
    output wire SUMA14_n;
    output wire SUMA15_n;
    output wire SUMA16_n;
    output wire SUMB13_n;
    output wire SUMB14_n;
    output wire SUMB15_n;
    output wire SUMB16_n;
    input wire US2SG;
    input wire WAG_n;
    input wire WALSG_n;
    input wire WBG_n;
    input wire WG1G_n;
    input wire WG2G_n;
    input wire WG3G_n;
    input wire WG4G_n;
    input wire WG5G_n;
    input wire WHOMPA;
    input wire WL01_n;
    input wire WL02_n;
    input wire WL12_n;
    output wire WL13;
    output wire WL13_n;
    output wire WL14;
    output wire WL14_n;
    output wire WL15;
    output wire WL15_n;
    output wire WL16;
    output wire WL16_n;
    input wire WLG_n;
    input wire WQG_n;
    input wire WYDG_n;
    input wire WYHIG_n;
    input wire WZG_n;
    input wire XUY01_n;
    input wire XUY02_n;
    output wire XUY13_n;
    output wire XUY14_n;
    inout wire Z15_n; //FPGA#wand
    inout wire Z16_n; //FPGA#wand
    wire __A11_1__X1;
    wire __A11_1__X1_n;
    wire __A11_1__X2;
    wire __A11_1__X2_n;
    wire __A11_1__Y1;
    wire __A11_1__Y1_n;
    wire __A11_1__Y2;
    wire __A11_1__Y2_n;
    wire __A11_1___A1_n;
    wire __A11_1___A2_n;
    wire __A11_1___B1_n;
    wire __A11_1___B2_n;
    wire __A11_1___CI_INTERNAL;
    wire __A11_1___Q1_n;
    wire __A11_1___Q2_n;
    wire __A11_1___RL_OUT_1;
    wire __A11_1___RL_OUT_2;
    wire __A11_1___Z1_n; //FPGA#wand
    wire __A11_1___Z2_n; //FPGA#wand
    wire __A11_2__X1;
    wire __A11_2__X1_n;
    wire __A11_2__X2;
    wire __A11_2__X2_n;
    wire __A11_2__Y1;
    wire __A11_2__Y1_n;
    wire __A11_2__Y2;
    wire __A11_2__Y2_n;
    wire __A11_2___B1_n;
    wire __A11_2___B2_n;
    wire __A11_2___CI_INTERNAL;
    wire __A11_2___CO_OUT; //FPGA#wand
    wire __A11_2___GEM1;
    wire __A11_2___Q1_n;
    wire __A11_2___Q2_n;
    wire __A11_2___RL_OUT_1;
    wire __A11_NET_130;
    wire __A11_NET_131;
    wire __A11_NET_132;
    wire __A11_NET_133;
    wire __A11_NET_134;
    wire __A11_NET_135;
    wire __A11_NET_136;
    wire __A11_NET_137;
    wire __A11_NET_138;
    wire __A11_NET_139;
    wire __A11_NET_140;
    wire __A11_NET_141;
    wire __A11_NET_142;
    wire __A11_NET_146;
    wire __A11_NET_147;
    wire __A11_NET_148;
    wire __A11_NET_149;
    wire __A11_NET_150;
    wire __A11_NET_151;
    wire __A11_NET_152;
    wire __A11_NET_154;
    wire __A11_NET_155;
    wire __A11_NET_156;
    wire __A11_NET_157;
    wire __A11_NET_160;
    wire __A11_NET_165;
    wire __A11_NET_166;
    wire __A11_NET_167;
    wire __A11_NET_168;
    wire __A11_NET_169;
    wire __A11_NET_170;
    wire __A11_NET_171;
    wire __A11_NET_172;
    wire __A11_NET_173;
    wire __A11_NET_174;
    wire __A11_NET_175;
    wire __A11_NET_176;
    wire __A11_NET_177;
    wire __A11_NET_178;
    wire __A11_NET_179;
    wire __A11_NET_180;
    wire __A11_NET_181;
    wire __A11_NET_182;
    wire __A11_NET_183;
    wire __A11_NET_184;
    wire __A11_NET_185;
    wire __A11_NET_186;
    wire __A11_NET_187;
    wire __A11_NET_188;
    wire __A11_NET_189;
    wire __A11_NET_190;
    wire __A11_NET_191;
    wire __A11_NET_192;
    wire __A11_NET_197;
    wire __A11_NET_198;
    wire __A11_NET_199;
    wire __A11_NET_200;
    wire __A11_NET_202;
    wire __A11_NET_203;
    wire __A11_NET_206;
    wire __A11_NET_207;
    wire __A11_NET_208;
    wire __A11_NET_209;
    wire __A11_NET_210;
    wire __A11_NET_211;
    wire __A11_NET_212;
    wire __A11_NET_213;
    wire __A11_NET_214;
    wire __A11_NET_215;
    wire __A11_NET_216;
    wire __A11_NET_217;
    wire __A11_NET_218;
    wire __A11_NET_219;
    wire __A11_NET_220;
    wire __A11_NET_221;
    wire __A11_NET_222;
    wire __A11_NET_223;
    wire __A11_NET_224;
    wire __A11_NET_225;
    wire __A11_NET_226;
    wire __A11_NET_227;
    wire __A11_NET_228;
    wire __A11_NET_229;
    wire __A11_NET_230;
    wire __A11_NET_231;
    wire __A11_NET_232;
    wire __A11_NET_233;
    wire __A11_NET_234;
    wire __A11_NET_235;
    wire __A11_NET_239;
    wire __A11_NET_240;
    wire __A11_NET_241;
    wire __A11_NET_242;
    wire __A11_NET_243;
    wire __A11_NET_244;
    wire __A11_NET_245;
    wire __A11_NET_247;
    wire __A11_NET_248;
    wire __A11_NET_249;
    wire __A11_NET_250;
    wire __A11_NET_253;
    wire __A11_NET_259;
    wire __A11_NET_260;
    wire __A11_NET_261;
    wire __A11_NET_262;
    wire __A11_NET_263;
    wire __A11_NET_264;
    wire __A11_NET_265;
    wire __A11_NET_266;
    wire __A11_NET_267;
    wire __A11_NET_268;
    wire __A11_NET_269;
    wire __A11_NET_270;
    wire __A11_NET_271;
    wire __A11_NET_272;
    wire __A11_NET_273;
    wire __A11_NET_274;
    wire __A11_NET_275;
    wire __A11_NET_276;
    wire __A11_NET_277;
    wire __A11_NET_278;
    wire __A11_NET_279;
    wire __A11_NET_280;
    wire __A11_NET_281;
    wire __A11_NET_282;
    wire __A11_NET_283;
    wire __A11_NET_284;
    wire __A11_NET_285;
    wire __A11_NET_286;
    wire __A11_NET_290;
    wire __A11_NET_291;
    wire __A11_NET_292;
    wire __A11_NET_293;
    wire __A11_NET_295;
    wire __A11_NET_296;
    wire __A11_NET_299;
    wire __A11_NET_300;
    wire __A11_NET_301;
    wire __A11_NET_302;
    wire __A11_NET_303;
    wire __A11_NET_304;
    wire __A11_NET_305;
    wire __A11_NET_306;
    wire __A11_NET_307;
    wire __A11_NET_308;
    wire __A11_NET_309;
    wire __A11_NET_310;
    wire __A11_NET_311;
    wire __A11_NET_312;
    wire __A11_NET_313;
    wire __A11_NET_314;
    wire __A11_NET_315;
    wire __CI15_n;
    wire __CO16; //FPGA#wand
    wire __G16_n; //FPGA#wand
    wire __L13_n; //FPGA#wand
    wire __L14_n; //FPGA#wand
    wire __RL16;
    wire __XUY15_n;
    wire __XUY16_n;

    pullup R11001(__CO16);
    pullup R11002(RL13_n);
    pullup R11003(__L13_n);
    pullup R11005(__A11_1___Z1_n);
    pullup R11006(G13_n);
    pullup R11007(RL14_n);
    pullup R11008(__L14_n);
    pullup R11009(__A11_1___Z2_n);
    pullup R11010(G14_n);
    pullup R11011(__A11_2___CO_OUT);
    pullup R11012(RL15_n);
    pullup R11013(L15_n);
    pullup R11015(Z15_n);
    pullup R11016(G15_n);
    pullup R11017(RL16_n);
    pullup R11018(L16_n);
    pullup R11019(Z16_n);
    pullup R11020(__G16_n);
    U74HC02 U11001(__A11_NET_197, A2XG_n, __A11_1___A1_n, __A11_NET_198, WYHIG_n, WL13_n, GND, WL12_n, WYDG_n, __A11_NET_192, __A11_1__Y1_n, CUG, __A11_1__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11002(MONEX, __A11_NET_197, __A11_1__X1_n, CLXC, CUG, __A11_1__X1, GND, __A11_1__Y1_n, __A11_NET_198, __A11_NET_192, __A11_1__Y1, __A11_1__X1_n, __A11_1__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11003(__A11_NET_202, __A11_1__X1_n, __A11_1__Y1_n, XUY13_n, __A11_1__X1, __A11_1__Y1, GND, __A11_NET_202, XUY13_n, __A11_NET_200, __A11_NET_202, SUMA13_n, __A11_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11004(__A11_NET_268, __A11_NET_270, SUMA13_n, SUMB13_n, RULOG_n, __A11_NET_180, GND, __A11_NET_184, __XUY15_n, XUY13_n, CI13_n, __A11_NET_271, __A11_NET_253, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U11005(CI13_n, __A11_NET_199, G13_n, GEM13, RL13_n, WL13, GND, WL13_n, WL13, MWL13, RL13_n, __A11_NET_146, __A11_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11006(SUMB13_n, __A11_NET_200, __A11_NET_199, __A11_NET_183, WAG_n, WL13_n, GND, WL15_n, WALSG_n, __A11_NET_185, __A11_1___A1_n, CAG, __A11_NET_181, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11007(__A11_NET_184, __CO16, __A11_NET_179, RL13_n, __A11_NET_188, __L13_n, GND, __A11_1___Z1_n, __A11_NET_214, RL13_n, __A11_NET_213, RL13_n, __A11_NET_215, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U11008(__A11_NET_178, RAG_n, __A11_1___A1_n, __A11_NET_182, WLG_n, WL13_n, GND, WL01_n, WALSG_n, __A11_NET_190, __L13_n, CLG2G, __A11_NET_191, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11009(__A11_NET_267, WG2G_n, WL16_n, __A11_NET_187, WQG_n, WL13_n, GND, __A11_NET_187, __A11_NET_186, __A11_1___Q1_n, __A11_1___Q1_n, CQG, __A11_NET_186, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11010(__A11_NET_189, RQG_n, __A11_1___Q1_n, __A11_NET_216, WZG_n, WL13_n, GND, __A11_NET_216, __A11_NET_217, __A11_NET_214, __A11_1___Z1_n, CZG, __A11_NET_217, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11011(__A11_1___RL_OUT_1, __A11_NET_189, MDT13, R1C, GND, __A11_NET_215, GND, __A11_NET_220, __A11_NET_219, __A11_NET_218, __A11_NET_203, __A11_NET_213, __A11_NET_212, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11012(__A11_NET_212, RZG_n, __A11_1___Z1_n, __A11_NET_221, WBG_n, WL13_n, GND, __A11_NET_221, __A11_NET_222, __A11_1___B1_n, __A11_1___B1_n, CBG, __A11_NET_222, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11013(__A11_NET_165, __CO16, __A11_NET_220, RL13_n, __A11_NET_208, G13_n, GND, G13_n, __A11_NET_211, RL14_n, __A11_NET_134, __L14_n, __A11_NET_137, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U11014(__A11_NET_219, RBHG_n, __A11_1___B1_n, __A11_NET_218, __A11_NET_222, RCG_n, GND, WL12_n, WG3G_n, __A11_NET_207, WL14_n, WG4G_n, __A11_NET_206, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11015(__A11_NET_183, __A11_NET_185, __A11_NET_180, __A11_NET_178, CH13, __A11_NET_179, GND, __A11_NET_188, __A11_NET_182, __A11_NET_190, __A11_NET_191, __A11_1___A1_n, __A11_NET_181, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11016(__A11_NET_210, L2GDG_n, L12_n, __A11_NET_209, WG1G_n, WL13_n, GND, G13_n, CGG, G13, RGG_n, G13_n, __A11_NET_203, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U11017(__A11_NET_210, __A11_NET_209, GND, __XUY16_n, XUY14_n, __A11_NET_165, GND, __A11_1___RL_OUT_1, RLG_n, __L13_n, GND, __A11_NET_211, G13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U11018(__A11_NET_208, GND, SA13, __A11_NET_207, __A11_NET_206,  , GND,  , GND, SA14, __A11_NET_157, __A11_NET_156, __A11_NET_155, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11019(__A11_NET_150, A2XG_n, __A11_1___A2_n, __A11_NET_154, WYHIG_n, WL14_n, GND, WL13_n, WYDG_n, __A11_NET_152, __A11_1__Y2_n, CUG, __A11_1__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11020(MONEX, __A11_NET_150, __A11_1__X2_n, CLXC, CUG, __A11_1__X2, GND, __A11_1__Y2_n, __A11_NET_154, __A11_NET_152, __A11_1__Y2, __A11_1__X2_n, __A11_1__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11021(__A11_NET_148, __A11_1__X2_n, __A11_1__Y2_n, XUY14_n, __A11_1__X2, __A11_1__Y2, GND, __G16_n, CGG, G16, __A11_NET_148, XUY14_n, __A11_NET_142, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U11022(__A11_NET_265, __A11_NET_267, __A11_NET_148, SUMA14_n, CO14, __CI15_n, GND, __A11_NET_147, SUMA14_n, SUMB14_n, RULOG_n, __A11_NET_266, G16, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11023(SUMB14_n, __A11_NET_142, __A11_NET_146, __A11_NET_149, WAG_n, WL14_n, GND, WL16_n, WALSG_n, __A11_NET_151, __A11_1___A2_n, CAG, __A11_NET_133, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11024(__A11_NET_149, __A11_NET_151, __A11_NET_147, __A11_NET_132, CH14, __A11_NET_134, GND, __A11_NET_137, __A11_NET_167, __A11_NET_166, __A11_NET_170, __A11_1___A2_n, __A11_NET_133, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11025(__A11_NET_132, RAG_n, __A11_1___A2_n, __A11_NET_167, WLG_n, WL14_n, GND, WL02_n, WALSG_n, __A11_NET_166, __L14_n, CLG2G, __A11_NET_170, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11026(RLG_n, __L14_n, __A11_1___RL_OUT_2, __A11_NET_135, __A11_NET_140, __A11_NET_136, GND, __A11_NET_131, MDT14, R1C, GND, __A11_1___RL_OUT_2, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11027(__A11_NET_169, WQG_n, WL14_n, __A11_1___Q2_n, __A11_NET_169, __A11_NET_139, GND, __A11_1___Q2_n, CQG, __A11_NET_139, RQG_n, __A11_1___Q2_n, __A11_NET_135, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11028(__A11_NET_136, RL14_n, __A11_NET_130, __A11_1___Z2_n, __A11_NET_131, RL14_n, GND, RL14_n, __A11_NET_177, G14_n, __A11_NET_155, G14_n, __A11_NET_171, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11029(__A11_NET_138, WZG_n, WL14_n, __A11_NET_130, __A11_NET_138, __A11_NET_141, GND, __A11_1___Z2_n, CZG, __A11_NET_141, RZG_n, __A11_1___Z2_n, __A11_NET_140, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11030(__A11_NET_168, WBG_n, WL14_n, __A11_1___B2_n, __A11_NET_168, __A11_NET_174, GND, __A11_1___B2_n, CBG, __A11_NET_174, RBHG_n, __A11_1___B2_n, __A11_NET_175, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U11031(__A11_NET_175, __A11_NET_176, __A11_NET_173, __A11_NET_172, G14, __A11_NET_171, GND, __A11_NET_259, GND, XUY02_n, __XUY16_n, __A11_NET_177, __A11_NET_160, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11032(__A11_NET_176, __A11_NET_174, RCG_n, __A11_NET_157, WL13_n, WG3G_n, GND, WL16_n, WG4G_n, __A11_NET_156, L2GDG_n, __L13_n, __A11_NET_173, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11033(__A11_NET_172, WG1G_n, WL14_n, G14, G14_n, CGG, GND, RGG_n, G14_n, __A11_NET_160, RGG_n, __G16_n, __A11_NET_253, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U11034(G14_n, GEM14, RL14_n, WL14, WL14, WL14_n, GND, MWL14, RL14_n,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11035(__A11_NET_290, A2XG_n, A15_n, __A11_NET_291, WYHIG_n, WL15_n, GND, WL14_n, WYDG_n, __A11_NET_286, __A11_2__Y1_n, CUG, __A11_2__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11036(BXVX, __A11_NET_290, __A11_2__X1_n, CLXC, CUG, __A11_2__X1, GND, __A11_2__Y1_n, __A11_NET_291, __A11_NET_286, __A11_2__Y1, __A11_2__X1_n, __A11_2__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11037(__A11_NET_295, __A11_2__X1_n, __A11_2__Y1_n, __XUY15_n, __A11_2__X1, __A11_2__Y1, GND, __A11_NET_295, __XUY15_n, __A11_NET_292, __A11_NET_295, SUMA15_n, __A11_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U11038(__A11_NET_303, __A11_NET_302, SUMA15_n, SUMB15_n, RULOG_n, __A11_NET_274, GND, __A11_NET_278, XUY01_n, __XUY15_n, __CI15_n, __A11_NET_304, G15, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U11039(__CI15_n, __A11_NET_293, G15_n, __A11_2___GEM1, RL15_n, WL15, GND, WL15_n, WL15, MWL15, RL15_n, __A11_NET_239, __A11_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11040(SUMB15_n, __A11_NET_292, __A11_NET_293, __A11_NET_277, WAG_n, WL15_n, GND, G16SW_n, WALSG_n, __A11_NET_279, A15_n, CAG, __A11_NET_275, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11041(__A11_NET_278, __A11_2___CO_OUT, __A11_NET_273, RL15_n, __A11_NET_282, L15_n, GND, Z15_n, __A11_NET_306, RL15_n, __A11_NET_307, RL15_n, __A11_NET_308, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 #(1'b1, 1'b0, 1'b1) U11042(__A11_NET_277, __A11_NET_279, __A11_NET_274, __A11_NET_272, CH16, __A11_NET_273, GND, __A11_NET_282, __A11_NET_276, __A11_NET_284, __A11_NET_285, A15_n, __A11_NET_275, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11043(__A11_NET_272, RAG_n, A15_n, __A11_NET_276, WLG_n, WL15_n, GND, G01_n, G2LSG_n, __A11_NET_284, L15_n, CLG1G, __A11_NET_285, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11044(__A11_NET_241, SUMA16_n, SUMA16_n, SUMB16_n, RUG_n, __A11_NET_240, GND, __A11_2___RL_OUT_1, RLG_n, L15_n, p4VSW, EAC_n, __CO16, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11045( ,  ,  , __A11_NET_281, WQG_n, WL15_n, GND, __A11_NET_281, __A11_NET_280, __A11_2___Q1_n, __A11_2___Q1_n, CQG, __A11_NET_280, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11046(__A11_NET_283, RQG_n, __A11_2___Q1_n, __A11_NET_309, WZG_n, WL15_n, GND, __A11_NET_309, __A11_NET_310, __A11_NET_306, Z15_n, CZG, __A11_NET_310, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11047(__A11_NET_305, RZG_n, Z15_n, __A11_NET_315, WBG_n, WL15_n, GND, __A11_NET_315, __A11_NET_314, __A11_2___B1_n, __A11_2___B1_n, CBG, __A11_NET_314, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11048(__A11_NET_312, RBHG_n, __A11_2___B1_n, __A11_NET_311, __A11_NET_314, RCG_n, GND, GND, p4VSW, __A11_NET_300, GND, p4VSW, __A11_NET_299, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11049(__A11_2___RL_OUT_1, __A11_NET_283, MDT15, R1C, __RL16, __A11_NET_308, GND, __A11_NET_313, __A11_NET_312, __A11_NET_311, __A11_NET_296, __A11_NET_307, __A11_NET_305, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11050(__A11_NET_259, __A11_2___CO_OUT, __A11_NET_313, RL15_n, __A11_NET_301, G15_n, GND, G15_n, __A11_NET_304, RL16_n, __A11_NET_227, L16_n, __A11_NET_228, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U11051(__A11_NET_303, L2GDG_n, __L14_n, __A11_NET_302, WG1G_n, WL15_n, GND, G15_n, CGG, G15, RGG_n, G15_n, __A11_NET_296, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U11052(__A11_NET_301, GND, SA16, __A11_NET_300, __A11_NET_299,  , GND,  , GND, SA16, __A11_NET_250, __A11_NET_249, __A11_NET_248, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11053(__A11_NET_243, A2XG_n, A16_n, __A11_NET_247, WYHIG_n, WL16_n, GND, WL16_n, WYDG_n, __A11_NET_245, __A11_2__Y2_n, CUG, __A11_2__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11054(MONEX, __A11_NET_243, __A11_2__X2_n, CLXC, CUG, __A11_2__X2, GND, __A11_2__Y2_n, __A11_NET_247, __A11_NET_245, __A11_2__Y2, __A11_2__X2_n, __A11_2__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11055(__A11_NET_241, __A11_2__X2_n, __A11_2__Y2_n, __XUY16_n, __A11_2__X2, __A11_2__Y2, GND,  ,  ,  , __A11_NET_241, __XUY16_n, __A11_NET_235, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11056(SUMB16_n, __A11_NET_235, __A11_NET_239, __A11_NET_242, WAG_n, WL16_n, GND, G16SW_n, WALSG_n, __A11_NET_244, A16_n, CAG, __A11_NET_226, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11057(__A11_NET_242, __A11_NET_244, __A11_NET_240, __A11_NET_225, CH16, __A11_NET_227, GND, __A11_NET_228, __A11_NET_263, __A11_NET_260, __A11_NET_264, A16_n, __A11_NET_226, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11058(__A11_NET_225, RAG_n, A16_n, __A11_NET_263, WLG_n, WL16_n, GND, __G16_n, G2LSG_n, __A11_NET_260, L16_n, CLG1G, __A11_NET_264, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11059(RLG_n, L16_n, __RL16, __A11_NET_230, __A11_NET_233, __A11_NET_229, GND, __A11_NET_223, MDT16, R1C, US2SG, __RL16, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11060(__A11_NET_262, WQG_n, WL16_n, __A11_2___Q2_n, __A11_NET_262, __A11_NET_232, GND, __A11_2___Q2_n, CQG, __A11_NET_232, RQG_n, __A11_2___Q2_n, __A11_NET_230, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11061(__A11_NET_229, RL16_n, __A11_NET_224, Z16_n, __A11_NET_223, RL16_n, GND, RL16_n, __A11_NET_271, __G16_n, __A11_NET_248, __G16_n, __A11_NET_266, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11062(__A11_NET_231, WZG_n, WL16_n, __A11_NET_224, __A11_NET_231, __A11_NET_234, GND, Z16_n, CZG, __A11_NET_234, RZG_n, Z16_n, __A11_NET_233, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11063(__A11_NET_261, WBG_n, WL16_n, __A11_2___B2_n, __A11_NET_261, __A11_NET_269, GND, __A11_2___B2_n, CBG, __A11_NET_269, RBHG_n, __A11_2___B2_n, __A11_NET_268, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11064(__A11_NET_270, __A11_NET_269, RCG_n, __A11_NET_250, WL14_n, WG3G_n, GND, WL01_n, WG5G_n, __A11_NET_249, L2GDG_n, L16_n, __A11_NET_265, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U11065(__G16_n, GEM16, RL16_n, WL16, WL16, WL16_n, GND, MWL16, RL16_n,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U11066(SUMA13_n, __A11_NET_202, XUY13_n, CI13_n, GND,  , GND,  , __A11_NET_148, XUY14_n, __A11_1___CI_INTERNAL, GND, SUMA14_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U11067(SUMA15_n, __A11_NET_295, __XUY15_n, __CI15_n, GND,  , GND,  , __A11_NET_241, __XUY16_n, __A11_2___CI_INTERNAL, WHOMPA, SUMA16_n, p4VSW, SIM_RST, SIM_CLK);
endmodule