`timescale 1ns/1ps
`default_nettype none

module inout_ii(VCC, GND, SIM_RST, SIM_CLK, GOJAM, F04B, FS05_n, F05A_n, F05B_n, TPOR_n, CCHG_n, WCHG_n, IN3301, ULLTHR, RRPONA, SMSEPR, RRRLSC, SPSRDY, ZEROP, S4BSAB, OPMSW2, LFTOFF, OPMSW3, GUIREL, STRPRS, OPCDFL, LVDAGD, IN3008, LRRLSC, IMUOPR, CH3310, CTLSAT, LEMATT, IMUCAG, IN3212, CDUFAL, HOLFUN, IN3213, IMUFAL, FREFUN, IN3214, ISSTOR, GCAPCL, IN3216, TEMPIN, TRST9, TRST10, PCHGOF, ROLGOF, MANpP, MANmP, MANpY, MANmY, MANpR, MANmR, TRANpX, TRANmX, TRANpY, TRANmY, TRANpZ, TRANmZ, MNIMpP, MNIMmP, MNIMpY, MNIMmY, MNIMpR, MNIMmR, PIPAFL, AGCWAR, OSCALM, CHWL01_n, CHWL02_n, CHWL03_n, CHWL04_n, CHWL05_n, CHWL06_n, CHWL07_n, CHWL08_n, CHWL09_n, CHWL10_n, CHWL11_n, CHWL12_n, CHWL13_n, CHWL14_n, CHWL16_n, CH1213, CH1214, CH1301, CH1302, CH1303, CH1304, CH1305, CH1306, CH1307, CH1308, CH1309, CH1310, CH1311, CH1316, CH1401, CH1402, CH1403, CH1404, CH1405, CH1406, CH1407, CH1408, CH1409, CH1410, CH1411, CH1412, CH1413, CH1414, CH1416, CH3312, XB0_n, XB1_n, XB2_n, XB3_n, XT1_n, XT3_n, WCH13_n, CCH11, RCH11_n, RCH33_n, WCH11_n, HNDRPT, CH3201, CH3202, CH3203, CH3204, CH3205, CH3206, CH3207, CH3208, CH3209, CH3210, CH3313, CH3314, CH3316, CHOR01_n, CHOR02_n, CHOR03_n, CHOR04_n, CHOR05_n, CHOR06_n, CHOR07_n, CHOR08_n, CHOR09_n, CHOR10_n, CHOR11_n, CHOR12_n, CHOR13_n, CHOR14_n, CHOR16_n);
    input wire VCC;
    input wire GND;
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire AGCWAR;
    output wire CCH11;
    input wire CCHG_n;
    input wire CDUFAL;
    input wire CH1213;
    input wire CH1214;
    input wire CH1301;
    input wire CH1302;
    input wire CH1303;
    input wire CH1304;
    input wire CH1305;
    input wire CH1306;
    input wire CH1307;
    input wire CH1308;
    input wire CH1309;
    input wire CH1310;
    input wire CH1311;
    input wire CH1316;
    input wire CH1401;
    input wire CH1402;
    input wire CH1403;
    input wire CH1404;
    input wire CH1405;
    input wire CH1406;
    input wire CH1407;
    input wire CH1408;
    input wire CH1409;
    input wire CH1410;
    input wire CH1411;
    input wire CH1412;
    input wire CH1413;
    input wire CH1414;
    input wire CH1416;
    output wire CH3201;
    output wire CH3202;
    output wire CH3203;
    output wire CH3204;
    output wire CH3205;
    output wire CH3206;
    output wire CH3207;
    output wire CH3208;
    output wire CH3209;
    output wire CH3210;
    input wire CH3310;
    input wire CH3312;
    output wire CH3313;
    output wire CH3314;
    output wire CH3316;
    output wire CHOR01_n; //FPGA#wand
    output wire CHOR02_n; //FPGA#wand
    output wire CHOR03_n; //FPGA#wand
    output wire CHOR04_n; //FPGA#wand
    output wire CHOR05_n; //FPGA#wand
    output wire CHOR06_n; //FPGA#wand
    output wire CHOR07_n; //FPGA#wand
    output wire CHOR08_n; //FPGA#wand
    output wire CHOR09_n; //FPGA#wand
    output wire CHOR10_n; //FPGA#wand
    output wire CHOR11_n; //FPGA#wand
    output wire CHOR12_n; //FPGA#wand
    output wire CHOR13_n; //FPGA#wand
    output wire CHOR14_n; //FPGA#wand
    output wire CHOR16_n; //FPGA#wand
    input wire CHWL01_n;
    input wire CHWL02_n;
    input wire CHWL03_n;
    input wire CHWL04_n;
    input wire CHWL05_n;
    input wire CHWL06_n;
    input wire CHWL07_n;
    input wire CHWL08_n;
    input wire CHWL09_n;
    input wire CHWL10_n;
    input wire CHWL11_n;
    input wire CHWL12_n;
    input wire CHWL13_n;
    input wire CHWL14_n;
    input wire CHWL16_n;
    input wire CTLSAT;
    input wire F04B;
    input wire F05A_n;
    input wire F05B_n;
    input wire FREFUN;
    input wire FS05_n;
    input wire GCAPCL;
    input wire GOJAM;
    input wire GUIREL;
    output wire HNDRPT;
    input wire HOLFUN;
    input wire IMUCAG;
    input wire IMUFAL;
    input wire IMUOPR;
    input wire IN3008;
    input wire IN3212;
    input wire IN3213;
    input wire IN3214;
    input wire IN3216;
    input wire IN3301;
    input wire ISSTOR;
    input wire LEMATT;
    input wire LFTOFF;
    input wire LRRLSC;
    input wire LVDAGD;
    input wire MANmP;
    input wire MANmR;
    input wire MANmY;
    input wire MANpP;
    input wire MANpR;
    input wire MANpY;
    input wire MNIMmP;
    input wire MNIMmR;
    input wire MNIMmY;
    input wire MNIMpP;
    input wire MNIMpR;
    input wire MNIMpY;
    input wire OPCDFL;
    input wire OPMSW2;
    input wire OPMSW3;
    input wire OSCALM;
    input wire PCHGOF;
    input wire PIPAFL;
    output wire RCH11_n;
    output wire RCH33_n;
    input wire ROLGOF;
    input wire RRPONA;
    input wire RRRLSC;
    input wire S4BSAB;
    input wire SMSEPR;
    input wire SPSRDY;
    input wire STRPRS;
    input wire TEMPIN;
    input wire TPOR_n;
    input wire TRANmX;
    input wire TRANmY;
    input wire TRANmZ;
    input wire TRANpX;
    input wire TRANpY;
    input wire TRANpZ;
    input wire TRST10;
    input wire TRST9;
    input wire ULLTHR;
    output wire WCH11_n;
    input wire WCH13_n;
    input wire WCHG_n;
    input wire XB0_n;
    input wire XB1_n;
    input wire XB2_n;
    input wire XB3_n;
    input wire XT1_n;
    input wire XT3_n;
    input wire ZEROP;
    wire __A17_1__F04B_n;
    wire __A17_1__FO5D;
    wire __A17_1__RCH30_n;
    wire __A17_1__RCH31_n;
    wire __A17_1__RCH32_n;
    wire __A17_1__TRP31A;
    wire __A17_1__TRP31B;
    wire __A17_1__TRP32;
    wire __A17_2__CCH10;
    wire __A17_2__RCH10_n;
    wire __A17_2__RLYB01;
    wire __A17_2__RLYB02;
    wire __A17_2__RLYB03;
    wire __A17_2__RLYB04;
    wire __A17_2__RLYB05;
    wire __A17_2__RLYB06;
    wire __A17_2__RLYB07;
    wire __A17_2__RLYB08;
    wire __A17_2__RLYB09;
    wire __A17_2__RLYB10;
    wire __A17_2__RLYB11;
    wire __A17_2__RYWD12;
    wire __A17_2__RYWD13;
    wire __A17_2__RYWD14;
    wire __A17_2__RYWD16;
    wire __A17_2__WCH10_n;
    wire __A17_NET_175;
    wire __A17_NET_176;
    wire __A17_NET_177;
    wire __A17_NET_178;
    wire __A17_NET_179;
    wire __A17_NET_180;
    wire __A17_NET_181;
    wire __A17_NET_182;
    wire __A17_NET_183;
    wire __A17_NET_184;
    wire __A17_NET_185;
    wire __A17_NET_186;
    wire __A17_NET_187;
    wire __A17_NET_188;
    wire __A17_NET_189;
    wire __A17_NET_190;
    wire __A17_NET_192; //FPGA#wand
    wire __A17_NET_193;
    wire __A17_NET_194;
    wire __A17_NET_195;
    wire __A17_NET_196;
    wire __A17_NET_197;
    wire __A17_NET_198;
    wire __A17_NET_199;
    wire __A17_NET_200;
    wire __A17_NET_201;
    wire __A17_NET_202;
    wire __A17_NET_203;
    wire __A17_NET_204;
    wire __A17_NET_205;
    wire __A17_NET_206;
    wire __A17_NET_207;
    wire __A17_NET_208;
    wire __A17_NET_209;
    wire __A17_NET_210;
    wire __A17_NET_211;
    wire __A17_NET_212;
    wire __A17_NET_213;
    wire __A17_NET_214;
    wire __A17_NET_215;
    wire __A17_NET_216;
    wire __A17_NET_217;
    wire __A17_NET_218;
    wire __A17_NET_219;
    wire __A17_NET_220;
    wire __A17_NET_221;
    wire __A17_NET_222;
    wire __A17_NET_223;
    wire __A17_NET_224;
    wire __A17_NET_225;
    wire __A17_NET_226;
    wire __A17_NET_227;
    wire __A17_NET_228;
    wire __A17_NET_229;
    wire __A17_NET_230;
    wire __A17_NET_231;
    wire __A17_NET_232;
    wire __A17_NET_233;
    wire __A17_NET_234;
    wire __A17_NET_235;
    wire __A17_NET_236;
    wire __A17_NET_237;
    wire __A17_NET_238;
    wire __A17_NET_239; //FPGA#wand
    wire __A17_NET_240;
    wire __A17_NET_241;
    wire __A17_NET_242;
    wire __A17_NET_243;
    wire __A17_NET_244;
    wire __A17_NET_246;
    wire __A17_NET_247;
    wire __A17_NET_249;
    wire __A17_NET_250; //FPGA#wand
    wire __A17_NET_251;
    wire __A17_NET_252;
    wire __A17_NET_253;
    wire __A17_NET_254;
    wire __A17_NET_255;
    wire __A17_NET_256;
    wire __A17_NET_257;
    wire __A17_NET_258;
    wire __A17_NET_259;
    wire __A17_NET_260;
    wire __A17_NET_261;
    wire __A17_NET_262;
    wire __A17_NET_263;
    wire __A17_NET_265;
    wire __A17_NET_266;
    wire __A17_NET_267;
    wire __A17_NET_268;
    wire __A17_NET_269;
    wire __A17_NET_270;
    wire __A17_NET_271;
    wire __A17_NET_272;
    wire __A17_NET_273;
    wire __A17_NET_274;
    wire __A17_NET_275;
    wire __A17_NET_276;
    wire __A17_NET_277;
    wire __A17_NET_278;
    wire __A17_NET_279;
    wire __A17_NET_280;
    wire __A17_NET_281;
    wire __A17_NET_282;
    wire __A17_NET_283;
    wire __A17_NET_284;
    wire __A17_NET_285;
    wire __A17_NET_286;
    wire __A17_NET_287;
    wire __A17_NET_288;
    wire __A17_NET_289;
    wire __A17_NET_290;
    wire __A17_NET_291;
    wire __A17_NET_292;
    wire __A17_NET_293;
    wire __A17_NET_294;
    wire __A17_NET_295;
    wire __A17_NET_296;
    wire __A17_NET_297;
    wire __A17_NET_298;
    wire __A17_NET_299;
    wire __A17_NET_300;
    wire __A17_NET_301;
    wire __A17_NET_302;
    wire __A17_NET_303;
    wire __A17_NET_304;
    wire __A17_NET_305;
    wire __A17_NET_306;
    wire __A17_NET_307;
    wire __A17_NET_308;
    wire __A17_NET_309;
    wire __A17_NET_310;
    wire __A17_NET_311;
    wire __A17_NET_312;
    wire __A17_NET_313;
    wire __A17_NET_314;
    wire __A17_NET_315;
    wire __A17_NET_316;
    wire __A17_NET_317;
    wire __A17_NET_318;
    wire __A17_NET_319;
    wire __A17_NET_321;
    wire __A17_NET_322;
    wire __A17_NET_324;
    wire __A17_NET_325;
    wire __A17_NET_326;
    wire __A17_NET_327;
    wire __A17_NET_328;
    wire __A17_NET_329;
    wire __A17_NET_330;
    wire __A17_NET_331;
    wire __A17_NET_332;
    wire __A17_NET_333;
    wire __A17_NET_334;
    wire __A17_NET_335;
    wire __A17_NET_336;
    wire __A17_NET_337;
    wire __A17_NET_338;
    wire __A17_NET_339;
    wire __A17_NET_340;
    wire __A17_NET_341;
    wire __A17_NET_342;
    wire __A17_NET_343;
    wire __A17_NET_344;
    wire __A17_NET_345;
    wire __A17_NET_346;
    wire __A17_NET_348;
    wire __A17_NET_349;
    wire __A17_NET_350;
    wire __A17_NET_351;
    wire __A17_NET_352;
    wire __A17_NET_353;
    wire __A17_NET_354;
    wire __A17_NET_355;
    wire __A17_NET_356;

    pullup R17001(CHOR01_n);
    pullup R17002(CHOR02_n);
    pullup R17003(CHOR03_n);
    pullup R17004(CHOR04_n);
    pullup R17005(CHOR05_n);
    pullup R17006(CHOR06_n);
    pullup R17007(CHOR07_n);
    pullup R17008(CHOR08_n);
    pullup R17009(CHOR09_n);
    pullup R17010(CHOR10_n);
    pullup R17011(CHOR11_n);
    pullup R17012(CHOR12_n);
    pullup R17013(CHOR13_n);
    pullup R17014(CHOR14_n);
    pullup R17015(CHOR16_n);
    pullup R17016(__A17_NET_192);
    pullup R17017(__A17_NET_239);
    pullup R17018(__A17_NET_250);
    U74HC02 U17001(__A17_NET_211, IN3301, RCH33_n, __A17_NET_212, XB3_n, XT3_n, GND, ULLTHR, __A17_1__RCH30_n, __A17_NET_209, XB0_n, XT3_n, __A17_NET_236, VCC, SIM_RST, SIM_CLK);
    U74HC04 U17002(__A17_NET_212, RCH33_n, __A17_NET_236, __A17_1__RCH30_n, __A17_NET_210, __A17_1__RCH31_n, GND, __A17_1__RCH32_n, __A17_NET_200, __A17_1__F04B_n, F04B, __A17_2__RLYB01, __A17_NET_331, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U17004(__A17_NET_258, CHOR01_n, __A17_NET_257, CHOR02_n, __A17_NET_260, CHOR03_n, GND, CHOR04_n, __A17_NET_259, CHOR05_n, __A17_NET_253, CHOR06_n, __A17_NET_251, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U17005(__A17_NET_215, MANpP, __A17_1__RCH31_n, __A17_NET_210, XB1_n, XT3_n, GND, SMSEPR, __A17_1__RCH30_n, __A17_NET_213, RRPONA, RCH33_n, __A17_NET_214, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17006(__A17_NET_204, MANmP, __A17_1__RCH31_n, __A17_NET_203, RRRLSC, RCH33_n, GND, MANpY, __A17_1__RCH31_n, __A17_NET_201, SPSRDY, __A17_1__RCH30_n, __A17_NET_202, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17007(__A17_NET_211, __A17_NET_209, __A17_NET_214, __A17_NET_213, __A17_NET_204, __A17_NET_257, GND, __A17_NET_260, __A17_NET_203, __A17_NET_202, __A17_NET_201, __A17_NET_258, __A17_NET_215, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17008(__A17_NET_207, S4BSAB, __A17_1__RCH30_n, __A17_NET_208, ZEROP, RCH33_n, GND, MANmY, __A17_1__RCH31_n, __A17_NET_206, LFTOFF, __A17_1__RCH30_n, __A17_NET_226, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17009(__A17_NET_208, __A17_NET_207, __A17_NET_205, __A17_NET_226, __A17_NET_225, __A17_NET_253, GND, __A17_NET_251, __A17_NET_224, __A17_NET_223, __A17_NET_230, __A17_NET_259, __A17_NET_206, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17010(__A17_NET_205, OPMSW2, RCH33_n, __A17_NET_225, MANpR, __A17_1__RCH31_n, GND, GUIREL, __A17_1__RCH30_n, __A17_NET_223, OPMSW3, RCH33_n, __A17_NET_224, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17011(__A17_NET_230, MANmR, __A17_1__RCH31_n, __A17_NET_228, OPCDFL, __A17_1__RCH30_n, GND, STRPRS, RCH33_n, __A17_NET_229, TRANpX, __A17_1__RCH31_n, __A17_NET_227, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17012(__A17_NET_229, __A17_NET_228, __A17_NET_219, __A17_NET_218, __A17_NET_217, __A17_NET_256, GND, __A17_NET_254, __A17_NET_216, __A17_NET_222, __A17_NET_221, __A17_NET_252, __A17_NET_227, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U17013(__A17_NET_252, CHOR07_n, __A17_NET_256, CHOR08_n, __A17_NET_254, CHOR09_n, GND, CHOR10_n, __A17_NET_255, CHOR11_n, __A17_NET_267, CHOR12_n, __A17_NET_266, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U17014(__A17_NET_218, IN3008, __A17_1__RCH30_n, __A17_NET_219, LVDAGD, RCH33_n, GND, TRANmX, __A17_1__RCH31_n, __A17_NET_217, IMUOPR, __A17_1__RCH30_n, __A17_NET_222, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17015(__A17_NET_216, LRRLSC, RCH33_n, __A17_NET_221, TRANpY, __A17_1__RCH31_n, GND, CTLSAT, __A17_1__RCH30_n, __A17_NET_220, TRANmY, __A17_1__RCH31_n, __A17_NET_185, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17016(CH3310, __A17_NET_220, __A17_NET_184, __A17_NET_183, __A17_NET_182, __A17_NET_267, GND, __A17_NET_266, __A17_NET_190, __A17_NET_189, __A17_NET_188, __A17_NET_255, __A17_NET_185, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17017(__A17_NET_183, IMUCAG, __A17_1__RCH30_n, __A17_NET_184, LEMATT, __A17_1__RCH32_n, GND, TRANpZ, __A17_1__RCH31_n, __A17_NET_182, CDUFAL, __A17_1__RCH30_n, __A17_NET_189, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17018(__A17_NET_190, IN3212, __A17_1__RCH32_n, __A17_NET_188, TRANmZ, __A17_1__RCH31_n, GND, IMUFAL, __A17_1__RCH30_n, __A17_NET_186, IN3213, __A17_1__RCH32_n, __A17_NET_187, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17019(__A17_NET_187, __A17_NET_186, __A17_NET_175, __A17_NET_176, __A17_NET_181, __A17_NET_268, GND, __A17_NET_269, __A17_NET_180, __A17_NET_178, __A17_NET_179, __A17_NET_270, __A17_NET_177, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U17020(__A17_NET_270, CHOR13_n, __A17_NET_268, CHOR14_n, __A17_NET_269, CHOR16_n, GND, __A17_NET_192, __A17_NET_262, __A17_NET_192, __A17_NET_261, __A17_NET_239, __A17_NET_265, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U17021(__A17_NET_177, HOLFUN, __A17_1__RCH31_n, __A17_NET_176, ISSTOR, __A17_1__RCH30_n, GND, IN3214, __A17_1__RCH32_n, __A17_NET_175, FREFUN, __A17_1__RCH31_n, __A17_NET_181, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17022(__A17_NET_178, TEMPIN, __A17_1__RCH30_n, __A17_NET_180, IN3216, __A17_1__RCH32_n, GND, GCAPCL, __A17_1__RCH31_n, __A17_NET_179, XB2_n, XT3_n, __A17_NET_200, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17023(MANpP, MANmP, MANmY, MANpR, MANmR, __A17_NET_261, GND, __A17_NET_197, __A17_NET_198, __A17_NET_192, F05A_n, __A17_NET_262, MANpY, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U17024(__A17_NET_195, CHWL12_n, WCH13_n, __A17_NET_198, __A17_NET_195, __A17_NET_199, GND, __A17_NET_197, __A17_NET_196, __A17_NET_194, __A17_1__F04B_n, FS05_n, __A17_1__FO5D, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17025(__A17_NET_198, GOJAM, __A17_NET_194, __A17_NET_192, __A17_1__FO5D, __A17_NET_196, GND, __A17_NET_265, TRANpX, TRANmX, TRANpY, __A17_NET_199, __A17_1__TRP31A, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U17026(__A17_1__TRP31A, __A17_NET_194, F05B_n, __A17_NET_240, __A17_NET_242, __A17_NET_241, GND, CHWL13_n, WCH13_n, __A17_NET_193, __A17_NET_240, F05B_n, __A17_1__TRP31B, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17027(TRANmY, TRANpZ, __A17_NET_243, __A17_NET_239, F05A_n, __A17_NET_242, GND, __A17_NET_241, __A17_NET_240, __A17_NET_239, __A17_1__FO5D, __A17_NET_263, TRANmZ, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U17028(__A17_NET_263, __A17_NET_239, __A17_NET_249, __A17_NET_250, __A17_NET_247, __A17_NET_250, GND, __A17_NET_250, __A17_NET_246, CHOR01_n, __A17_NET_327, CHOR07_n, __A17_NET_341, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 U17029(__A17_NET_243, GOJAM, MNIMpR, MNIMmR, TRST9, __A17_NET_247, GND, __A17_NET_246, TRST10, PCHGOF, ROLGOF, __A17_NET_244, __A17_1__TRP31B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17030(__A17_NET_243, __A17_NET_193, __A17_NET_244, CH3201, MNIMpP, __A17_1__RCH32_n, GND, MNIMmP, __A17_1__RCH32_n, CH3202, MNIMpY, __A17_1__RCH32_n, CH3203, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17031(CH3204, MNIMmY, __A17_1__RCH32_n, CH3205, MNIMpR, __A17_1__RCH32_n, GND, MNIMmR, __A17_1__RCH32_n, CH3206, TRST9, __A17_1__RCH32_n, CH3207, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U17032(CH3208, TRST10, __A17_1__RCH32_n, CH3209, PCHGOF, __A17_1__RCH32_n, GND, ROLGOF, __A17_1__RCH32_n, CH3210, __A17_NET_235, __A17_NET_234, __A17_NET_233, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U17033(__A17_NET_249, MNIMpP, MNIMmP, MNIMpY, MNIMmY,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U17034(WCHG_n, XT1_n, __A17_NET_237, __A17_NET_250, F05A_n, __A17_NET_235, GND, __A17_NET_234, __A17_NET_233, __A17_1__FO5D, __A17_NET_250, __A17_NET_297, XB1_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U17035(__A17_1__TRP32, __A17_NET_233, F05B_n, __A17_NET_232, CHWL14_n, WCH13_n, GND, __A17_NET_232, __A17_NET_231, __A17_NET_237, __A17_NET_238, TPOR_n, HNDRPT, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17036(__A17_NET_237, GOJAM, __A17_1__TRP31A, __A17_1__TRP31B, __A17_1__TRP32, __A17_NET_238, GND, __A17_NET_327, CH1301, __A17_NET_326, CH1401, __A17_NET_231, __A17_1__TRP32, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17037(CH3313, PIPAFL, RCH33_n, CH3314, AGCWAR, RCH33_n, GND, OSCALM, RCH33_n, CH3316, CHWL01_n, __A17_2__WCH10_n, __A17_NET_329, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17038(__A17_NET_331, __A17_NET_329, __A17_NET_330, __A17_NET_330, __A17_NET_331, __A17_2__CCH10, GND, __A17_NET_331, __A17_2__RCH10_n, __A17_NET_326, CHWL02_n, __A17_2__WCH10_n, __A17_NET_328, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17039(__A17_NET_335, __A17_NET_328, __A17_NET_334, __A17_NET_334, __A17_NET_335, __A17_2__CCH10, GND, __A17_NET_335, __A17_2__RCH10_n, __A17_NET_333, CHWL03_n, __A17_2__WCH10_n, __A17_NET_316, VCC, SIM_RST, SIM_CLK);
    U74HC04 U17040(__A17_NET_335, __A17_2__RLYB02, __A17_NET_317, __A17_2__RLYB03, __A17_NET_324, __A17_2__RLYB04, GND, __A17_2__RLYB05, __A17_NET_321, __A17_2__RLYB06, __A17_NET_354, __A17_2__RLYB07, __A17_NET_353, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17041(CH1302, __A17_NET_333, CH1303, __A17_NET_312, CH1403, __A17_NET_311, GND, __A17_NET_318, CH1304, __A17_NET_325, CH1404, __A17_NET_332, CH1402, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U17042(__A17_NET_332, CHOR02_n, __A17_NET_311, CHOR03_n, __A17_NET_318, CHOR04_n, GND, CHOR05_n, __A17_NET_348, CHOR06_n, __A17_NET_356, CHOR08_n, __A17_NET_345, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17043(__A17_NET_317, __A17_NET_316, __A17_NET_315, __A17_NET_315, __A17_NET_317, __A17_2__CCH10, GND, __A17_NET_317, __A17_2__RCH10_n, __A17_NET_312, CHWL04_n, __A17_2__WCH10_n, __A17_NET_313, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17044(__A17_NET_324, __A17_NET_313, __A17_NET_314, __A17_NET_314, __A17_NET_324, __A17_2__CCH10, GND, __A17_NET_324, __A17_2__RCH10_n, __A17_NET_325, CHWL05_n, __A17_2__WCH10_n, __A17_NET_322, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17045(__A17_NET_321, __A17_NET_322, __A17_NET_319, __A17_NET_319, __A17_NET_321, __A17_2__CCH10, GND, __A17_NET_321, __A17_2__RCH10_n, __A17_NET_350, CHWL06_n, __A17_2__WCH10_n, __A17_NET_346, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17046(CH1305, __A17_NET_350, CH1306, __A17_NET_355, CH1406, __A17_NET_356, GND,  ,  ,  ,  , __A17_NET_348, CH1405, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17047(__A17_NET_354, __A17_NET_346, __A17_NET_349, __A17_NET_349, __A17_NET_354, __A17_2__CCH10, GND, __A17_NET_354, __A17_2__RCH10_n, __A17_NET_355, CHWL07_n, __A17_2__WCH10_n, __A17_NET_351, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17048(__A17_NET_353, __A17_NET_351, __A17_NET_352, __A17_NET_352, __A17_NET_353, __A17_2__CCH10, GND, __A17_NET_353, __A17_2__RCH10_n, __A17_NET_340, CHWL08_n, __A17_2__WCH10_n, __A17_NET_336, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17049(CH1307, __A17_NET_340, CH1308, __A17_NET_339, CH1408, __A17_NET_345, GND, __A17_NET_288, CH1309, __A17_NET_287, CH1409, __A17_NET_341, CH1407, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17050(__A17_NET_338, __A17_NET_336, __A17_NET_337, __A17_NET_337, __A17_NET_338, __A17_2__CCH10, GND, __A17_NET_338, __A17_2__RCH10_n, __A17_NET_339, CHWL09_n, __A17_2__WCH10_n, __A17_NET_344, VCC, SIM_RST, SIM_CLK);
    U74HC04 U17051(__A17_NET_338, __A17_2__RLYB08, __A17_NET_343, __A17_2__RLYB09, __A17_NET_285, __A17_2__RLYB10, GND, __A17_2__RLYB11, __A17_NET_291, __A17_2__RYWD12, __A17_NET_272, __A17_2__RYWD13, __A17_NET_281, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17052(__A17_NET_343, __A17_NET_344, __A17_NET_342, __A17_NET_342, __A17_NET_343, __A17_2__CCH10, GND, __A17_NET_343, __A17_2__RCH10_n, __A17_NET_287, CHWL10_n, __A17_2__WCH10_n, __A17_NET_284, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U17053(__A17_NET_288, CHOR09_n, __A17_NET_292, CHOR10_n, __A17_NET_274, CHOR11_n, GND, CHOR12_n, __A17_NET_273, CHOR13_n, __A17_NET_279, CHOR14_n, __A17_NET_301, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17054(__A17_NET_285, __A17_NET_284, __A17_NET_283, __A17_NET_283, __A17_NET_285, __A17_2__CCH10, GND, __A17_NET_285, __A17_2__RCH10_n, __A17_NET_286, CHWL11_n, __A17_2__WCH10_n, __A17_NET_290, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17055(CH1310, __A17_NET_286, CH1311, __A17_NET_275, CH1411, __A17_NET_274, GND, __A17_NET_273, CH3312, __A17_NET_271, CH1412, __A17_NET_292, CH1410, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17056(__A17_NET_291, __A17_NET_290, __A17_NET_289, __A17_NET_289, __A17_NET_291, __A17_2__CCH10, GND, __A17_NET_291, __A17_2__RCH10_n, __A17_NET_275, CHWL12_n, __A17_2__WCH10_n, __A17_NET_277, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17057(__A17_NET_272, __A17_NET_277, __A17_NET_276, __A17_NET_276, __A17_NET_272, __A17_2__CCH10, GND, __A17_NET_272, __A17_2__RCH10_n, __A17_NET_271, CHWL13_n, __A17_2__WCH10_n, __A17_NET_280, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17058(__A17_NET_281, __A17_NET_280, __A17_NET_282, __A17_NET_282, __A17_NET_281, __A17_2__CCH10, GND, __A17_NET_281, __A17_2__RCH10_n, __A17_NET_278, CHWL14_n, __A17_2__WCH10_n, __A17_NET_303, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17059(__A17_NET_305, __A17_NET_303, __A17_NET_304, __A17_NET_304, __A17_NET_305, __A17_2__CCH10, GND, __A17_NET_305, __A17_2__RCH10_n, __A17_NET_302, CHWL16_n, __A17_2__WCH10_n, __A17_NET_309, VCC, SIM_RST, SIM_CLK);
    U74HC04 U17060(__A17_NET_305, __A17_2__RYWD14, __A17_NET_308, __A17_2__RYWD16, __A17_NET_296, __A17_2__WCH10_n, GND, __A17_2__CCH10, __A17_NET_295, WCH11_n, __A17_NET_297, CCH11, __A17_NET_298, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17061(__A17_NET_308, __A17_NET_309, __A17_NET_310, __A17_NET_310, __A17_NET_308, __A17_2__CCH10, GND, __A17_NET_308, __A17_2__RCH10_n, __A17_NET_306, __A17_NET_294, GOJAM, __A17_NET_295, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U17062(__A17_NET_307, CHOR16_n,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK); //FPGA#OD:2
    U74HC27 U17063(CH1213, __A17_NET_278, CH1214, __A17_NET_302, CH1414, __A17_NET_301, GND, __A17_NET_307, CH1316, __A17_NET_306, CH1416, __A17_NET_279, CH1413, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17064(WCHG_n, XB0_n, CCHG_n, XT1_n, XB0_n, __A17_NET_294, GND, __A17_NET_299, CCHG_n, XT1_n, XB1_n, __A17_NET_296, XT1_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17065(__A17_NET_293, XT1_n, XB0_n, __A17_NET_298, __A17_NET_299, GOJAM, GND, XT1_n, XB1_n, __A17_NET_300,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U17066(__A17_NET_293, __A17_2__RCH10_n, __A17_NET_300, RCH11_n,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
endmodule