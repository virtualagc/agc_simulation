`include "components/agc_parts.v"

module timer(VCC, GND, SIM_RST, CLOCK, MSTRTP, MSTP, PHS2, PHS2_n, PHS3_n, PHS4, PHS4_n, RT, RT_n, WT, WT_n, CT, CT_n, CLK, TT_n, P01, P01_n, P02, P02_n, P03, P03_n, P04, P04_n, P05, P05_n, SBY, ALGA, STRT1, STRT2, GOJ1, STOPA, GOJAM, GOJAM_n, STOP, STOP_n, WL15, WL15_n, WL16, WL16_n, FS01_n, T01, T01_n, T02, T02_n, T03, T03_n, T04, T04_n, T05, T05_n, T06, T06_n, T07, T07_n, T08, T08_n, T09, T09_n, T10, T10_n, T11, T11_n, T12, T12_n, OVF_n, UNF_n, MONWT, Q2A, MGOJAM, MSTPIT_n);
    input wire SIM_RST;
    input wire ALGA;
    output wire CLK;
    input wire CLOCK;
    output wire CT;
    output wire CT_n;
    output wire FS01_n;
    input wire GND;
    input wire GOJ1;
    output wire GOJAM;
    output wire GOJAM_n;
    output wire MGOJAM;
    output wire MONWT;
    input wire MSTP;
    output wire MSTPIT_n;
    input wire MSTRTP;
    wire NET_117;
    wire NET_131;
    wire NET_132;
    wire NET_133;
    wire NET_134;
    wire NET_135;
    wire NET_136;
    wire NET_137;
    wire NET_138;
    wire NET_139;
    wire NET_140;
    wire NET_141;
    wire NET_142;
    wire NET_143;
    wire NET_144;
    wire NET_145;
    wire NET_146;
    wire NET_147;
    wire NET_148;
    wire NET_149;
    wire NET_150;
    wire NET_151;
    wire NET_152;
    wire NET_153;
    wire NET_154;
    wire NET_155;
    wire NET_156;
    wire NET_157;
    wire NET_158;
    wire NET_159;
    wire NET_160;
    wire NET_161;
    wire NET_162;
    wire NET_163;
    wire NET_164;
    wire NET_165;
    wire NET_166;
    wire NET_167;
    wire NET_168;
    wire NET_169;
    wire NET_170;
    wire NET_171;
    wire NET_172;
    wire NET_173;
    wire NET_174;
    wire NET_175;
    wire NET_176;
    wire NET_177;
    wire NET_178;
    wire NET_179;
    wire NET_180;
    wire NET_181;
    wire NET_182;
    output wire OVF_n;
    output wire P01;
    output wire P01_n;
    output wire P02;
    output wire P02_n;
    output wire P03;
    output wire P03_n;
    output wire P04;
    output wire P04_n;
    output wire P05;
    output wire P05_n;
    output wire PHS2;
    output wire PHS2_n;
    output wire PHS3_n;
    output wire PHS4;
    output wire PHS4_n;
    output wire Q2A;
    output wire RT;
    output wire RT_n;
    input wire SBY;
    output wire STOP;
    output wire STOPA;
    output wire STOP_n;
    input wire STRT1;
    input wire STRT2;
    output wire T01;
    output wire T01_n;
    output wire T02;
    output wire T02_n;
    output wire T03;
    output wire T03_n;
    output wire T04;
    output wire T04_n;
    output wire T05;
    output wire T05_n;
    output wire T06;
    output wire T06_n;
    output wire T07;
    output wire T07_n;
    output wire T08;
    output wire T08_n;
    output wire T09;
    output wire T09_n;
    output wire T10;
    output wire T10_n;
    output wire T11;
    output wire T11_n;
    output wire T12;
    output wire T12_n;
    output wire TT_n;
    output wire UNF_n;
    input wire VCC;
    input wire WL15;
    input wire WL15_n;
    input wire WL16;
    input wire WL16_n;
    output wire WT;
    output wire WT_n;
    wire __A02_1__EVNSET_n;
    wire __A02_1__ODDSET_n;
    wire __A02_1__OVFSTB_n;
    wire __A02_1__RINGA_n;
    wire __A02_1__RINGB_n;
    wire __A02_1__cdiv_1__A;
    wire __A02_1__cdiv_1__B;
    wire __A02_1__cdiv_1__D;
    wire __A02_1__cdiv_1__FS;
    wire __A02_1__cdiv_1__FS_n;
    wire __A02_1__cdiv_2__A;
    wire __A02_1__cdiv_2__B;
    wire __A02_1__cdiv_2__C;
    wire __A02_1__cdiv_2__D;
    wire __A02_1__cdiv_2__F;
    wire __A02_1__cdiv_2__FS;
    wire __A02_1__cdiv_2__FS_n;
    wire __A02_1__evnset;
    wire __A02_1__oddset;
    wire __A02_1__ovfstb_r1;
    wire __A02_1__ovfstb_r2;
    wire __A02_1__ovfstb_r3;
    wire __A02_1__ovfstb_r4;
    wire __A02_1__ovfstb_r5;
    wire __A02_1__ovfstb_r6;
    wire __A02_2__F01A;
    wire __A02_2__F01B;
    wire __A02_2__F01C;
    wire __A02_2__F01D;
    wire __A02_2__FS01;
    wire __A02_3__MT01;
    wire __A02_3__MT02;
    wire __A02_3__MT03;
    wire __A02_3__MT04;
    wire __A02_3__MT05;
    wire __A02_3__MT06;
    wire __A02_3__MT07;
    wire __A02_3__MT08;
    wire __A02_3__MT09;
    wire __A02_3__MT10;
    wire __A02_3__MT11;
    wire __A02_3__MT12;
    wire __A02_3__OVF;
    wire __A02_3__T01DC_n;
    wire __A02_3__T02DC_n;
    wire __A02_3__T03DC_n;
    wire __A02_3__T04DC_n;
    wire __A02_3__T05DC_n;
    wire __A02_3__T06DC_n;
    wire __A02_3__T07DC_n;
    wire __A02_3__T08DC_n;
    wire __A02_3__T09DC_n;
    wire __A02_3__T10DC_n;
    wire __A02_3__T12DC_n;
    wire __A02_3__T12SET;
    wire __A02_3__UNF;

    pullup R2001(NET_142);
    pullup R2002(__A02_3__T12SET);
    U74HC02 #(0, 1, 0, 0) U2001(__A02_1__cdiv_1__D, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__B, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__B, __A02_1__cdiv_1__FS, GND, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__A, __A02_1__cdiv_1__FS, __A02_1__cdiv_1__A, __A02_1__cdiv_1__FS, PHS2, VCC, SIM_RST);
    wire U2002_8_NC;
    wire U2002_9_NC;
    wire U2002_10_NC;
    wire U2002_11_NC;
    U74HC27 #(0, 1, 0) U2002(__A02_1__cdiv_1__D, CLOCK, __A02_1__cdiv_1__B, CLOCK, PHS2, __A02_1__cdiv_1__A, GND, U2002_8_NC, U2002_9_NC, U2002_10_NC, U2002_11_NC, __A02_1__cdiv_1__B, __A02_1__cdiv_1__A, VCC, SIM_RST);
    U74HC04 #(1, 0, 0, 1, 0, 0) U2003(__A02_1__cdiv_1__D, __A02_1__cdiv_2__F, PHS2, PHS2_n, PHS4, PHS4_n, GND, NET_117, __A02_1__cdiv_1__B, CT, NET_117, CT_n, CT, VCC, SIM_RST);
    wire U2004_8_NC;
    wire U2004_9_NC;
    wire U2004_10_NC;
    wire U2004_11_NC;
    wire U2004_12_NC;
    wire U2004_13_NC;
    U74HC02 U2004(PHS4, __A02_1__cdiv_2__F, __A02_1__cdiv_1__A, __A02_1__oddset, STOP, __A02_1__RINGA_n, GND, U2004_8_NC, U2004_9_NC, U2004_10_NC, U2004_11_NC, U2004_12_NC, U2004_13_NC, VCC, SIM_RST);
    U74HC04 U2005(__A02_1__cdiv_1__FS_n, WT, WT, WT_n, WT, TT_n, GND, __A02_1__ovfstb_r5, __A02_1__ovfstb_r4, __A02_1__ovfstb_r6, __A02_1__ovfstb_r5, __A02_1__OVFSTB_n, __A02_1__ovfstb_r2, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U2006(__A02_1__cdiv_2__D, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__FS, GND, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__A, __A02_1__cdiv_2__FS, __A02_1__cdiv_2__A, __A02_1__cdiv_2__FS, __A02_1__cdiv_2__C, VCC, SIM_RST);
    wire U2007_8_NC;
    wire U2007_9_NC;
    wire U2007_10_NC;
    wire U2007_11_NC;
    U74HC27 #(0, 1, 0) U2007(__A02_1__cdiv_2__D, __A02_1__cdiv_2__F, __A02_1__cdiv_2__B, __A02_1__cdiv_2__F, __A02_1__cdiv_2__C, __A02_1__cdiv_2__A, GND, U2007_8_NC, U2007_9_NC, U2007_10_NC, U2007_11_NC, __A02_1__cdiv_2__B, __A02_1__cdiv_2__A, VCC, SIM_RST);
    U74HC04 #(1, 0, 1, 0, 0, 0) U2008(__A02_1__cdiv_2__D, __A02_1__RINGA_n, __A02_1__oddset, __A02_1__ODDSET_n, __A02_1__cdiv_2__C, __A02_1__RINGB_n, GND, __A02_1__evnset, __A02_1__RINGB_n, __A02_1__EVNSET_n, __A02_1__evnset, RT, __A02_1__cdiv_1__A, VCC, SIM_RST);
    U74HC02 U2009(__A02_1__ovfstb_r1, CT_n, __A02_1__ovfstb_r2, __A02_1__ovfstb_r2, __A02_1__ovfstb_r6, __A02_1__ovfstb_r1, GND, __A02_1__ovfstb_r4, __A02_1__ovfstb_r2, __A02_1__ovfstb_r3, __A02_1__ovfstb_r3, __A02_1__ovfstb_r1, __A02_1__ovfstb_r4, VCC, SIM_RST);
    wire U2010_12_NC;
    wire U2010_13_NC;
    U74HC04 #(1, 0, 0, 0, 0, 0) U2010(CT, PHS3_n, WT_n, CLK, WT_n, MONWT, GND, Q2A, WT_n, RT_n, RT, U2010_12_NC, U2010_13_NC, VCC, SIM_RST);
    U74HC27 U2011(__A02_1__RINGB_n, P05_n, P04, P05, __A02_1__RINGA_n, NET_152, GND, NET_145, GND, NET_142, __A02_1__EVNSET_n, NET_151, P04_n, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U2012(P01, NET_151, P01_n, P01_n, P01, NET_152, GND, __A02_1__RINGA_n, P01, NET_148, P01_n, __A02_1__RINGB_n, NET_153, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U2013(P02, NET_148, P02_n, P02_n, P02, NET_153, GND, __A02_1__RINGB_n, P02, NET_150, P02_n, __A02_1__RINGA_n, NET_149, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U2014(P03, NET_150, P03_n, P03_n, P03, NET_149, GND, __A02_1__RINGA_n, P03, NET_135, P03_n, __A02_1__RINGB_n, NET_136, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U2015(P04, NET_135, P04_n, P04_n, P04, NET_136, GND, __A02_1__RINGB_n, P04, NET_138, P04_n, __A02_1__RINGA_n, NET_137, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U2016(P05, NET_138, P05_n, P05_n, P05, NET_137, GND, NET_142, GOJ1, NET_134, __A02_1__EVNSET_n, NET_133, NET_146, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U2017(__A02_2__F01D, FS01_n, __A02_2__F01B, FS01_n, __A02_2__F01B, __A02_2__FS01, GND, FS01_n, __A02_2__F01A, __A02_2__FS01, __A02_2__F01A, __A02_2__FS01, __A02_2__F01C, VCC, SIM_RST);
    wire U2018_8_NC;
    wire U2018_9_NC;
    wire U2018_10_NC;
    wire U2018_11_NC;
    U74HC27 #(0, 1, 0) U2018(__A02_2__F01D, P01_n, __A02_2__F01B, P01_n, __A02_2__F01C, __A02_2__F01A, GND, U2018_8_NC, U2018_9_NC, U2018_10_NC, U2018_11_NC, __A02_2__F01B, __A02_2__F01A, VCC, SIM_RST);
    U74HC27 #(1, 1, 0) U2019(SBY, ALGA, STRT1, STRT2, NET_134, NET_132, GND, NET_140, GND, NET_141, __A02_1__EVNSET_n, NET_131, MSTRTP, VCC, SIM_RST);
    wire U2020_5_NC;
    wire U2020_6_NC;
    wire U2020_8_NC;
    wire U2020_9_NC;
    wire U2020_10_NC;
    wire U2020_11_NC;
    wire U2020_12_NC;
    wire U2020_13_NC;
    U74LVC07 U2020(NET_131, NET_142, NET_132, NET_142, U2020_5_NC, U2020_6_NC, GND, U2020_8_NC, U2020_9_NC, U2020_10_NC, U2020_11_NC, U2020_12_NC, U2020_13_NC, VCC, SIM_RST);
    U74HC04 #(1, 0, 1, 0, 1, 0) U2021(NET_142, NET_133, MSTP, NET_141, GOJAM_n, GOJAM, GND, MGOJAM, GOJAM, STOP, STOP_n, MSTPIT_n, STOP, VCC, SIM_RST);
    wire U2022_11_NC;
    wire U2022_12_NC;
    wire U2022_13_NC;
    U74HC02 U2022(NET_139, __A02_1__EVNSET_n, MSTP, GOJAM_n, STRT2, STOPA, GND, STOPA, NET_143, STOP_n, U2022_11_NC, U2022_12_NC, U2022_13_NC, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 1) U2023(NET_144, NET_145, STOPA, STOPA, NET_144, NET_146, GND, NET_140, NET_143, NET_147, NET_147, NET_139, NET_143, VCC, SIM_RST);
    U74HC27 #(1, 0, 0) U2024(__A02_3__T12SET, GOJAM, __A02_3__T01DC_n, NET_177, GOJAM, NET_174, GND, NET_177, __A02_3__T02DC_n, NET_175, GOJAM, __A02_3__T12DC_n, NET_176, VCC, SIM_RST);
    U74HC02 #(0, 0, 0, 1) U2025(NET_176, __A02_3__T12DC_n, NET_174, NET_164, __A02_3__T12DC_n, __A02_1__ODDSET_n, GND, __A02_3__T12DC_n, __A02_1__EVNSET_n, T12, NET_164, NET_174, __A02_3__T01DC_n, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U2026(NET_169, __A02_3__T01DC_n, __A02_1__EVNSET_n, T01, __A02_3__T01DC_n, __A02_1__ODDSET_n, GND, NET_169, NET_177, __A02_3__T02DC_n, __A02_3__T02DC_n, __A02_1__ODDSET_n, NET_168, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U2027(T02, __A02_3__T02DC_n, __A02_1__EVNSET_n, __A02_3__T03DC_n, NET_168, NET_175, GND, __A02_3__T03DC_n, __A02_1__EVNSET_n, NET_170, __A02_3__T03DC_n, __A02_1__ODDSET_n, T03, VCC, SIM_RST);
    U74HC27 U2028(__A02_3__T03DC_n, NET_171, __A02_3__T04DC_n, NET_172, GOJAM, NET_171, GND, NET_172, __A02_3__T05DC_n, NET_173, GOJAM, NET_175, GOJAM, VCC, SIM_RST);
    U74HC02 #(1, 0, 0, 1) U2029(__A02_3__T04DC_n, NET_170, NET_171, NET_165, __A02_3__T04DC_n, __A02_1__ODDSET_n, GND, __A02_3__T04DC_n, __A02_1__EVNSET_n, T04, NET_165, NET_172, __A02_3__T05DC_n, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U2030(NET_155, __A02_3__T05DC_n, __A02_1__EVNSET_n, T05, __A02_3__T05DC_n, __A02_1__ODDSET_n, GND, NET_173, NET_155, __A02_3__T06DC_n, __A02_1__EVNSET_n, __A02_3__T06DC_n, T06, VCC, SIM_RST);
    U74HC27 U2031(GOJAM, NET_180, GOJAM, NET_179, __A02_3__T07DC_n, NET_180, GND, NET_179, GOJAM, NET_182, __A02_3__T08DC_n, NET_173, __A02_3__T06DC_n, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U2032(NET_167, __A02_1__ODDSET_n, __A02_3__T06DC_n, __A02_3__T07DC_n, NET_180, NET_167, GND, __A02_1__ODDSET_n, __A02_3__T07DC_n, T07, __A02_1__EVNSET_n, __A02_3__T07DC_n, NET_166, VCC, SIM_RST);
    U74HC02 #(1, 0, 0, 1) U2033(__A02_3__T08DC_n, NET_179, NET_166, T08, __A02_1__EVNSET_n, __A02_3__T08DC_n, GND, __A02_1__ODDSET_n, __A02_3__T08DC_n, NET_159, NET_182, NET_159, __A02_3__T09DC_n, VCC, SIM_RST);
    U74HC27 U2034(GOJAM, NET_181, GOJAM, NET_178, __A02_3__T10DC_n, NET_181, GND, NET_178, GOJAM, NET_160, NET_163, NET_182, __A02_3__T09DC_n, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U2035(T09, __A02_1__ODDSET_n, __A02_3__T09DC_n, NET_162, __A02_1__EVNSET_n, __A02_3__T09DC_n, GND, NET_181, NET_162, __A02_3__T10DC_n, __A02_1__EVNSET_n, NET_181, NET_160, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U2036(NET_161, __A02_1__ODDSET_n, __A02_3__T10DC_n, NET_163, NET_178, NET_161, GND, __A02_1__EVNSET_n, __A02_3__T10DC_n, T10, __A02_1__ODDSET_n, NET_163, T11, VCC, SIM_RST);
    wire U2037_4_NC;
    wire U2037_5_NC;
    wire U2037_6_NC;
    wire U2037_8_NC;
    wire U2037_9_NC;
    wire U2037_10_NC;
    wire U2037_11_NC;
    wire U2037_12_NC;
    wire U2037_13_NC;
    U74HC02 U2037(NET_154, NET_177, NET_174, U2037_4_NC, U2037_5_NC, U2037_6_NC, GND, U2037_8_NC, U2037_9_NC, U2037_10_NC, U2037_11_NC, U2037_12_NC, U2037_13_NC, VCC, SIM_RST);
    U74HC27 U2038(NET_172, NET_171, NET_182, NET_181, __A02_1__EVNSET_n, NET_158, GND, NET_157, NET_173, NET_180, NET_179, NET_156, NET_175, VCC, SIM_RST);
    wire U2039_10_NC;
    wire U2039_11_NC;
    wire U2039_12_NC;
    wire U2039_13_NC;
    U74LVC07 U2039(NET_154, __A02_3__T12SET, NET_156, __A02_3__T12SET, NET_158, __A02_3__T12SET, GND, __A02_3__T12SET, NET_157, U2039_10_NC, U2039_11_NC, U2039_12_NC, U2039_13_NC, VCC, SIM_RST);
    U74HC04 U2040(T01, T01_n, T01_n, __A02_3__MT01, T02, T02_n, GND, __A02_3__MT02, T02_n, T03_n, T03, __A02_3__MT03, T03_n, VCC, SIM_RST);
    U74HC04 U2041(T04, T04_n, T04_n, __A02_3__MT04, T05, T05_n, GND, __A02_3__MT05, T05_n, T06_n, T06, __A02_3__MT06, T06_n, VCC, SIM_RST);
    U74HC04 U2042(T07, T07_n, T07_n, __A02_3__MT07, T08, T08_n, GND, __A02_3__MT08, T08_n, T09_n, T09, __A02_3__MT09, T09_n, VCC, SIM_RST);
    U74HC04 U2043(T10, T10_n, T10_n, __A02_3__MT10, T11, T11_n, GND, __A02_3__MT11, T11_n, T12_n, T12, __A02_3__MT12, T12_n, VCC, SIM_RST);
    wire U2044_8_NC;
    wire U2044_9_NC;
    wire U2044_10_NC;
    wire U2044_11_NC;
    U74HC27 U2044(WL15_n, WL16, __A02_1__OVFSTB_n, WL15, WL16_n, __A02_3__UNF, GND, U2044_8_NC, U2044_9_NC, U2044_10_NC, U2044_11_NC, __A02_3__OVF, __A02_1__OVFSTB_n, VCC, SIM_RST);
    wire U2045_5_NC;
    wire U2045_6_NC;
    wire U2045_8_NC;
    wire U2045_9_NC;
    wire U2045_10_NC;
    wire U2045_11_NC;
    wire U2045_12_NC;
    wire U2045_13_NC;
    U74HC04 U2045(__A02_3__OVF, OVF_n, __A02_3__UNF, UNF_n, U2045_5_NC, U2045_6_NC, GND, U2045_8_NC, U2045_9_NC, U2045_10_NC, U2045_11_NC, U2045_12_NC, U2045_13_NC, VCC, SIM_RST);
endmodule