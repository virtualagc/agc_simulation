`timescale 1ns/1ps
`default_nettype none

module alarms(SIM_RST, SIM_CLK, p4VDC, p4VSW, GND, GOJAM, PHS2_n, PHS3_n, PHS4_n, T02_n, T03_n, T04_n, T07_n, T09_n, T10, T10_n, T11_n, T12_n, CT, CT_n, P02, P02_n, P03, P03_n, SB0_n, SB1_n, SB2_n, FS01, F05A_n, F05B_n, F07A, F07B_n, F08B, FS09, FS10, F10A_n, F10B, F12B, FS13, FS14, F14B, FS17, F17A, F17B, ST0_n, ST1_n, STRT2, VFAIL, n2FSFAL, FLTOUT, SCAFAL, SBY, STNDBY_n, CTROR, CTROR_n, PSEUDO, TC0, TCF0, GNHNC, NISQL_n, IIP, IIP_n, PALE, PIPAFL, TEMPIN, TMPOUT, CCH33, CA6_n, XB7_n, ALTEST, ERRST, DOSCAL, DBLTST, MSTRT, NHALGA, NHVFAL, MLOAD, MREAD, MLDCH, MRDCH, MNHNC, T1P, T2P, T3P, T4P, T5P, T6P, CDUXP, CDUXM, CDUYP, CDUYM, CDUZP, CDUZM, TRNP, TRNM, SHAFTP, SHAFTM, PIPXP, PIPXM, PIPYP, PIPYM, PIPZP, PIPZM, BMAGXP, BMAGXM, BMAGYP, BMAGYM, BMAGZP, BMAGZM, INLNKP, INLNKM, RNRADP, RNRADM, GYROD, CDUXD, CDUYD, CDUZD, TRUND, SHAFTD, THRSTD, EMSD, OTLNKM, ALTM, ALGA, STRT1, BKTF_n, RSSB, CHINC, CHINC_n, FETCH0, FETCH0_n, FETCH1, STORE1_n, STFET1_n, INCSET_n, INKL, INKL_n, INOTLD, MON_n, MONpCH, MSTRTP, AGCWAR, OSCALM, TMPCAU, RESTRT, MRPTAL_n, MTCAL_n, MCTRAL_n, MVFAIL_n, MWARNF_n, MSCAFL_n, MSCDBL_n, MOSCAL_n, MPIPAL_n, MWATCH_n, MINKL, MREQIN);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VDC;
    input wire p4VSW;
    input wire GND;
    output wire AGCWAR;
    output wire ALGA;
    input wire ALTEST;
    input wire ALTM;
    output wire BKTF_n;
    input wire BMAGXM;
    input wire BMAGXP;
    input wire BMAGYM;
    input wire BMAGYP;
    input wire BMAGZM;
    input wire BMAGZP;
    input wire CA6_n;
    input wire CCH33;
    input wire CDUXD;
    input wire CDUXM;
    input wire CDUXP;
    input wire CDUYD;
    input wire CDUYM;
    input wire CDUYP;
    input wire CDUZD;
    input wire CDUZM;
    input wire CDUZP;
    output wire CHINC;
    output wire CHINC_n;
    input wire CT;
    input wire CTROR;
    input wire CTROR_n;
    input wire CT_n;
    input wire DBLTST;
    input wire DOSCAL;
    input wire EMSD;
    input wire ERRST;
    input wire F05A_n;
    input wire F05B_n;
    input wire F07A;
    input wire F07B_n;
    input wire F08B;
    input wire F10A_n;
    input wire F10B;
    input wire F12B;
    input wire F14B;
    input wire F17A;
    input wire F17B;
    output wire FETCH0;
    output wire FETCH0_n;
    output wire FETCH1;
    input wire FLTOUT;
    input wire FS01;
    input wire FS09;
    input wire FS10;
    input wire FS13;
    input wire FS14;
    input wire FS17;
    input wire GNHNC;
    input wire GOJAM;
    input wire GYROD;
    input wire IIP;
    input wire IIP_n;
    output wire INCSET_n;
    output wire INKL;
    output wire INKL_n;
    input wire INLNKM;
    input wire INLNKP;
    output wire INOTLD;
    output wire MCTRAL_n; //FPGA#wand
    output wire MINKL; //FPGA#wand
    input wire MLDCH;
    input wire MLOAD;
    input wire MNHNC;
    output wire MON_n;
    output wire MONpCH;
    output wire MOSCAL_n; //FPGA#wand
    output wire MPIPAL_n; //FPGA#wand
    input wire MRDCH;
    input wire MREAD;
    output wire MREQIN; //FPGA#wand
    output wire MRPTAL_n; //FPGA#wand
    output wire MSCAFL_n; //FPGA#wand
    output wire MSCDBL_n; //FPGA#wand
    input wire MSTRT;
    output wire MSTRTP;
    output wire MTCAL_n; //FPGA#wand
    output wire MVFAIL_n; //FPGA#wand
    output wire MWARNF_n; //FPGA#wand
    output wire MWATCH_n; //FPGA#wand
    input wire NHALGA;
    input wire NHVFAL;
    input wire NISQL_n;
    output wire OSCALM;
    input wire OTLNKM;
    input wire P02;
    input wire P02_n;
    input wire P03;
    input wire P03_n;
    input wire PALE;
    input wire PHS2_n;
    input wire PHS3_n;
    input wire PHS4_n;
    input wire PIPAFL;
    input wire PIPXM;
    input wire PIPXP;
    input wire PIPYM;
    input wire PIPYP;
    input wire PIPZM;
    input wire PIPZP;
    input wire PSEUDO;
    output wire RESTRT;
    input wire RNRADM;
    input wire RNRADP;
    output wire RSSB;
    input wire SB0_n;
    input wire SB1_n;
    input wire SB2_n;
    input wire SBY;
    input wire SCAFAL;
    input wire SHAFTD;
    input wire SHAFTM;
    input wire SHAFTP;
    input wire ST0_n;
    input wire ST1_n;
    output wire STFET1_n;
    input wire STNDBY_n;
    output wire STORE1_n;
    output wire STRT1;
    input wire STRT2;
    input wire T02_n;
    input wire T03_n;
    input wire T04_n;
    input wire T07_n;
    input wire T09_n;
    input wire T10;
    input wire T10_n;
    input wire T11_n;
    input wire T12_n;
    input wire T1P;
    input wire T2P;
    input wire T3P;
    input wire T4P;
    input wire T5P;
    input wire T6P;
    input wire TC0;
    input wire TCF0;
    input wire TEMPIN;
    input wire THRSTD;
    output wire TMPCAU;
    input wire TMPOUT;
    input wire TRNM;
    input wire TRNP;
    input wire TRUND;
    input wire VFAIL;
    input wire XB7_n;
    wire __A13_1__CGCWAR;
    wire __A13_1__CKTAL_n; //FPGA#wand
    wire __A13_1__CON1;
    wire __A13_1__CON2;
    wire __A13_1__CON3;
    wire __A13_1__DOFILT;
    wire __A13_1__F12B_n;
    wire __A13_1__F14H;
    wire __A13_1__FILTIN;
    wire __A13_1__FS13_n;
    wire __A13_1__NOTEST;
    wire __A13_1__NOTEST_n;
    wire __A13_1__SBYEXT;
    wire __A13_1__SCADBL;
    wire __A13_1__SCAS10;
    wire __A13_1__SCAS17;
    wire __A13_1__SYNC14_n;
    wire __A13_1__SYNC4_n;
    wire __A13_1__TEMPIN_n;
    wire __A13_1__WARN;
    wire __A13_1__WATCH;
    wire __A13_1__WATCHP;
    wire __A13_2__INOTRD;
    wire __A13_2__STORE1;
    input wire n2FSFAL;
    wire net_R13002_Pad2; //FPGA#wand
    wire net_R13003_Pad2; //FPGA#wand
    wire net_R13004_Pad2; //FPGA#wand
    wire net_U13001_Pad13;
    wire net_U13001_Pad2;
    wire net_U13001_Pad6;
    wire net_U13001_Pad8;
    wire net_U13002_Pad1;
    wire net_U13002_Pad10;
    wire net_U13002_Pad12;
    wire net_U13003_Pad1;
    wire net_U13003_Pad10;
    wire net_U13003_Pad13;
    wire net_U13003_Pad3;
    wire net_U13004_Pad10;
    wire net_U13004_Pad4;
    wire net_U13004_Pad5;
    wire net_U13004_Pad6;
    wire net_U13004_Pad8;
    wire net_U13004_Pad9;
    wire net_U13005_Pad10;
    wire net_U13005_Pad11;
    wire net_U13005_Pad13;
    wire net_U13006_Pad11;
    wire net_U13006_Pad13;
    wire net_U13006_Pad5;
    wire net_U13006_Pad9;
    wire net_U13007_Pad10;
    wire net_U13007_Pad6;
    wire net_U13007_Pad8;
    wire net_U13008_Pad1;
    wire net_U13008_Pad11;
    wire net_U13008_Pad2;
    wire net_U13009_Pad13;
    wire net_U13010_Pad1;
    wire net_U13010_Pad10;
    wire net_U13011_Pad1;
    wire net_U13011_Pad13;
    wire net_U13012_Pad1;
    wire net_U13012_Pad10;
    wire net_U13012_Pad12;
    wire net_U13012_Pad13;
    wire net_U13012_Pad3;
    wire net_U13013_Pad10;
    wire net_U13013_Pad11;
    wire net_U13013_Pad12;
    wire net_U13013_Pad8;
    wire net_U13013_Pad9;
    wire net_U13014_Pad1;
    wire net_U13014_Pad3;
    wire net_U13029_Pad1;
    wire net_U13029_Pad10;
    wire net_U13029_Pad13;
    wire net_U13029_Pad2;
    wire net_U13029_Pad3;
    wire net_U13029_Pad8;
    wire net_U13030_Pad10;
    wire net_U13030_Pad4;
    wire net_U13030_Pad6;
    wire net_U13030_Pad8;
    wire net_U13031_Pad12;
    wire net_U13031_Pad13;
    wire net_U13031_Pad4;
    wire net_U13031_Pad8;
    wire net_U13031_Pad9;
    wire net_U13032_Pad12;
    wire net_U13034_Pad13;
    wire net_U13035_Pad1;
    wire net_U13035_Pad13;
    wire net_U13036_Pad11;
    wire net_U13037_Pad11;
    wire net_U13037_Pad12;
    wire net_U13037_Pad5;
    wire net_U13038_Pad1;
    wire net_U13038_Pad10;
    wire net_U13038_Pad13;
    wire net_U13039_Pad1;
    wire net_U13039_Pad13;
    wire net_U13039_Pad4;
    wire net_U13039_Pad9;
    wire net_U13040_Pad4;
    wire net_U13042_Pad13;
    wire net_U13042_Pad8;
    wire net_U13043_Pad13;
    wire net_U13044_Pad10;
    wire net_U13044_Pad8;
    wire net_U13044_Pad9;
    wire net_U13045_Pad1;
    wire net_U13052_Pad1;
    wire net_U13115_Pad10;
    wire net_U13115_Pad12;
    wire net_U13115_Pad13;
    wire net_U13115_Pad9;
    wire net_U13116_Pad10;
    wire net_U13116_Pad13;
    wire net_U13117_Pad8;
    wire net_U13118_Pad1;
    wire net_U13118_Pad10;
    wire net_U13119_Pad12;
    wire net_U13119_Pad6;
    wire net_U13119_Pad8;
    wire net_U13120_Pad10;
    wire net_U13120_Pad12;
    wire net_U13120_Pad13;
    wire net_U13122_Pad10;
    wire net_U13122_Pad13;
    wire net_U13123_Pad13;
    wire net_U13124_Pad4;
    wire net_U13125_Pad1;
    wire net_U13125_Pad10;
    wire net_U13125_Pad13;
    wire net_U13125_Pad3;
    wire net_U13125_Pad4;
    wire net_U13126_Pad6;
    wire net_U13127_Pad5;

    pullup R13001(__A13_1__CKTAL_n);
    pullup R13002(net_R13002_Pad2);
    pullup R13003(net_R13003_Pad2);
    pullup R13004(net_R13004_Pad2);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U13001(MSTRT, net_U13001_Pad2, F12B, __A13_1__F12B_n, __A13_1__F14H, net_U13001_Pad6, GND, net_U13001_Pad8, net_R13002_Pad2, __A13_1__NOTEST, __A13_1__NOTEST_n, __A13_1__DOFILT, net_U13001_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U13002(net_U13002_Pad1, F05B_n, net_U13001_Pad2, net_U13002_Pad12, net_U13002_Pad1, net_U13002_Pad10, GND, net_U13002_Pad12, net_U13001_Pad2, net_U13002_Pad10, F05A_n, net_U13002_Pad12, MSTRTP, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U13003(net_U13003_Pad1, IIP, net_U13003_Pad3, net_U13003_Pad3, net_U13003_Pad1, F14B, GND, IIP_n, net_U13003_Pad13, net_U13003_Pad10, net_U13003_Pad10, F14B, net_U13003_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U13004(__A13_1__F12B_n, FS14, PALE, net_U13004_Pad4, net_U13004_Pad5, net_U13004_Pad6, GND, net_U13004_Pad8, net_U13004_Pad9, net_U13004_Pad10, __A13_1__WATCHP, __A13_1__F14H, __A13_1__FS13_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U13005(net_U13004_Pad4, net_U13003_Pad3, net_U13001_Pad6, net_U13004_Pad5, net_U13003_Pad13, net_U13001_Pad6, GND, net_U13004_Pad4, net_U13004_Pad5, net_U13005_Pad10, net_U13005_Pad11, F10B, net_U13005_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U13006(net_U13004_Pad6, __A13_1__CKTAL_n, net_U13004_Pad8, __A13_1__CKTAL_n, net_U13006_Pad5, net_R13002_Pad2, GND, net_R13002_Pad2, net_U13006_Pad9, net_R13002_Pad2, net_U13006_Pad11, net_R13002_Pad2, net_U13006_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 #(1'b1, 1'b0, 1'b0) U13007(TC0, TCF0, T12_n, PHS4_n, NISQL_n, net_U13007_Pad6, GND, net_U13007_Pad8, __A13_1__NOTEST, net_U13007_Pad10, T09_n, net_U13005_Pad11, net_U13005_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U13008(net_U13008_Pad1, net_U13008_Pad2, net_U13008_Pad11, net_U13008_Pad11, net_U13008_Pad1, F10B, GND, net_U13005_Pad13, F10A_n, net_U13004_Pad9, net_U13008_Pad11, F10A_n, net_U13004_Pad10, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b0, 1'b1) U13009(net_U13008_Pad2, TCF0, TC0, INKL, T04_n,  , GND,  , INLNKP, INLNKM, RNRADP, RNRADM, net_U13009_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U13010(net_U13010_Pad1, net_U13004_Pad9, net_U13004_Pad10, net_U13007_Pad10, net_U13001_Pad8, net_U13010_Pad10, GND, net_U13007_Pad10, INKL, net_U13010_Pad10, PSEUDO, NISQL_n, __A13_1__NOTEST_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U13011(net_U13011_Pad1, GYROD, CDUXD, CDUYD, CDUZD,  , GND,  , TRUND, SHAFTD, THRSTD, EMSD, net_U13011_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U13012(net_U13012_Pad1, net_U13007_Pad8, net_U13012_Pad3, net_U13012_Pad3, net_U13012_Pad1, INKL, GND, T03_n, net_U13012_Pad1, net_U13012_Pad10, net_U13012_Pad10, net_U13012_Pad12, net_U13012_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U13013(INKL, T03_n, net_U13012_Pad10, net_U13012_Pad12, GOJAM, net_U13001_Pad13, GND, net_U13013_Pad8, net_U13013_Pad9, net_U13013_Pad10, net_U13013_Pad11, net_U13013_Pad12, CTROR, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U13014(net_U13014_Pad1, net_U13013_Pad12, net_U13014_Pad3, net_U13014_Pad3, net_U13014_Pad1, F07A, GND, net_U13014_Pad3, F07B_n, net_U13012_Pad12, NHALGA, __A13_1__CKTAL_n, ALGA, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U13115(__A13_1__SCAS10, __A13_1__CON2, FS10, __A13_1__SCAS17, FS17, DOSCAL, GND, F05B_n, net_U13115_Pad9, net_U13115_Pad10, net_U13115_Pad10, net_U13115_Pad12, net_U13115_Pad13, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U13116(VFAIL, net_U13115_Pad9,  ,  , TEMPIN, __A13_1__TEMPIN_n, GND,  ,  , net_U13116_Pad10, F14B, __A13_1__FILTIN, net_U13116_Pad13, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U13117(net_U13115_Pad13, net_U13115_Pad9, F05A_n, net_U13115_Pad13, NHVFAL, net_U13052_Pad1, GND, net_U13117_Pad8, F05A_n, net_U13115_Pad13, STNDBY_n, net_U13115_Pad12, NHVFAL, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U13118(net_U13118_Pad1, net_U13052_Pad1, STRT1, STRT1, net_U13118_Pad1, net_U13118_Pad10, GND, net_U13115_Pad12, F05A_n, net_U13118_Pad10, __A13_1__CON3, n2FSFAL, __A13_1__SCADBL, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U13119(net_U13117_Pad8, __A13_1__DOFILT, SB0_n, net_R13003_Pad2, net_U13116_Pad10, net_U13119_Pad6, GND, net_U13119_Pad8, FLTOUT, SCAFAL, AGCWAR, net_U13119_Pad12, __A13_1__SCADBL, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U13120(__A13_1__CON3, __A13_1__CON2, FS10,  ,  ,  , GND, ALTEST, net_U13120_Pad13, net_U13120_Pad10, net_R13003_Pad2, net_U13120_Pad12, net_U13120_Pad13, p4VDC, SIM_RST, SIM_CLK);
    U74LVC07 U13121(net_U13119_Pad12, net_R13003_Pad2, net_U13120_Pad10, net_R13003_Pad2,  ,  , GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK); //FPGA#OD:2,4
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U13122(net_U13120_Pad12, SB2_n, net_U13116_Pad10, net_U13116_Pad13, net_U13119_Pad6, net_U13122_Pad10, GND, net_U13116_Pad13, F08B, net_U13122_Pad10, FLTOUT, SCAFAL, net_U13122_Pad13, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U13123(net_U13122_Pad13, __A13_1__WARN, __A13_1__WARN, __A13_1__CGCWAR,  ,  , GND,  ,  ,  ,  , TMPCAU, net_U13123_Pad13, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U13124(AGCWAR, net_U13119_Pad8, CCH33, net_U13124_Pad4, STRT2, OSCALM, GND, net_U13124_Pad4, CCH33, OSCALM, __A13_1__TEMPIN_n, TMPOUT, net_U13123_Pad13, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U13125(net_U13125_Pad1, GOJAM, net_U13125_Pad3, net_U13125_Pad4, ALTEST, net_U13125_Pad3, GND, SBY, net_U13125_Pad13, net_U13125_Pad10, net_U13125_Pad10, T10, net_U13125_Pad13, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U13126(net_U13125_Pad1, ERRST, CT_n, P02_n, P03, net_U13126_Pad6, GND,  ,  ,  ,  , net_U13125_Pad3, __A13_1__SBYEXT, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U13127(net_U13125_Pad4, RESTRT, net_U13125_Pad10, __A13_1__SBYEXT, net_U13127_Pad5, __A13_1__SYNC4_n, GND, __A13_1__SYNC14_n, net_U13126_Pad6,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC4002 U13128(net_U13127_Pad5, FS01, P02, P03_n, CT_n,  , GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U13029(net_U13029_Pad1, net_U13029_Pad2, net_U13029_Pad3, net_U13029_Pad3, net_U13029_Pad1, F17B, GND, net_U13029_Pad8, SB1_n, net_U13029_Pad10, __A13_1__WATCHP, __A13_1__WATCH, net_U13029_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U13030(SB2_n, net_U13029_Pad3, net_U13013_Pad9, net_U13030_Pad4, net_U13013_Pad11, net_U13030_Pad6, GND, net_U13030_Pad8, net_U13013_Pad9, net_U13030_Pad10, net_U13013_Pad11, __A13_1__WATCHP, net_U13029_Pad8, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b1) U13031(__A13_1__WATCH, net_U13029_Pad13, net_U13029_Pad10, net_U13031_Pad4, OTLNKM, ALTM, GND, net_U13031_Pad8, net_U13031_Pad9, net_U13013_Pad11, net_U13013_Pad8, net_U13031_Pad12, net_U13031_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U13032( ,  , net_R13004_Pad2, net_U13013_Pad9, MLOAD, net_U13013_Pad10, GND, net_U13030_Pad4, MREAD, net_U13030_Pad10, MLDCH, net_U13032_Pad12, MRDCH, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U13033(net_U13006_Pad9, T5P, T6P, CDUXP, CDUXM,  , GND,  , CDUYP, CDUYM, CDUZP, CDUZM, net_U13006_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U13034(net_U13006_Pad13, TRNP, TRNM, SHAFTP, SHAFTM,  , GND,  , PIPXP, PIPXM, PIPYP, PIPYM, net_U13034_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U13035(net_U13035_Pad1, PIPZP, PIPZM, BMAGXP, BMAGXM,  , GND,  , BMAGYP, BMAGYM, BMAGZP, BMAGZM, net_U13035_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U13036(net_U13011_Pad1, net_R13002_Pad2, net_U13011_Pad13, net_R13002_Pad2, net_U13031_Pad4, net_R13002_Pad2, GND, net_R13004_Pad2, net_U13007_Pad6, net_R13004_Pad2, net_U13036_Pad11, net_R13002_Pad2, net_U13034_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 U13037(net_U13013_Pad9, net_U13032_Pad12, net_U13013_Pad11, GOJAM, net_U13037_Pad5, net_U13031_Pad9, GND, net_U13031_Pad12, net_U13031_Pad13, GOJAM, net_U13037_Pad11, net_U13037_Pad12, net_U13013_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U13038(net_U13038_Pad1, MRDCH, MLDCH, MREAD, MLOAD,  , GND,  , net_U13031_Pad12, net_U13038_Pad10, INOTLD, __A13_2__INOTRD, net_U13038_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b0, 1'b1) U13039(net_U13039_Pad1, net_U13030_Pad6, net_U13038_Pad10, net_U13039_Pad4, net_U13030_Pad8, INOTLD, GND, net_U13039_Pad4, net_U13039_Pad9, INOTLD, net_U13037_Pad12, __A13_2__INOTRD, net_U13039_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U13040(net_U13039_Pad1, GOJAM, MON_n, net_U13040_Pad4, ST1_n, net_U13037_Pad11, GND, net_U13039_Pad9, T12_n, CT, PHS2_n, net_U13038_Pad10, net_U13037_Pad11, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U13041(__A13_2__INOTRD, net_U13039_Pad13, net_U13039_Pad9, __A13_2__STORE1, ST1_n, net_U13031_Pad13, GND, ST1_n, net_U13039_Pad1, FETCH1, net_U13031_Pad12, net_U13038_Pad10, MON_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U13042(FETCH0, ST0_n, MON_n, STFET1_n, __A13_2__STORE1, FETCH1, GND, net_U13042_Pad8, T11_n, net_U13037_Pad5, CTROR_n, net_U13031_Pad9, net_U13042_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U13043(net_U13039_Pad9, net_U13040_Pad4, __A13_2__STORE1, STORE1_n, FETCH0, FETCH0_n, GND, MONpCH, net_U13038_Pad13,  ,  , INCSET_n, net_U13043_Pad13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U13044(FETCH1, __A13_2__STORE1, net_U13042_Pad13, T12_n, PHS3_n, net_U13044_Pad10, GND, net_U13044_Pad8, net_U13044_Pad9, net_U13044_Pad10, GOJAM, net_U13042_Pad8, CHINC, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b0, 1'b1) U13045(net_U13045_Pad1, net_U13013_Pad9, MNHNC, net_U13031_Pad9, CTROR_n,  , GND,  , T1P, T2P, T3P, T4P, net_U13006_Pad5, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U13046(net_U13044_Pad9, net_U13045_Pad1, net_U13044_Pad8, net_U13043_Pad13, T02_n, net_U13044_Pad9, GND, net_U13044_Pad8, MONpCH, INKL_n, __A13_2__INOTRD, INOTLD, CHINC_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U13047(INKL_n, INKL,  ,  , T10_n, BKTF_n, GND, CHINC, CHINC_n, __A13_1__FS13_n, FS13, __A13_1__CON1, DBLTST, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U13048(net_U13044_Pad9, T07_n, T02_n, CA6_n, XB7_n, net_U13029_Pad2, GND,  ,  ,  ,  , RSSB, PHS3_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U13049(net_U13036_Pad11, GNHNC, PSEUDO, net_U13031_Pad8, PHS2_n, net_U13038_Pad1, GND, __A13_1__CON1, FS09, __A13_1__CON2,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U13050( ,  ,  ,  ,  ,  , GND,  ,  ,  ,  , net_U13029_Pad8, F17A, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U13051(net_U13035_Pad1, net_R13002_Pad2, net_U13035_Pad13, net_R13002_Pad2, net_U13009_Pad13, net_R13002_Pad2, GND, MRPTAL_n, net_U13005_Pad10, MTCAL_n, net_U13010_Pad1, MCTRAL_n, net_U13012_Pad13, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74LVC06 U13052(net_U13052_Pad1, MVFAIL_n, PIPAFL, MPIPAL_n, __A13_1__SCADBL, MSCDBL_n, GND, MWATCH_n, __A13_1__WATCH, MSCAFL_n, SCAFAL, MWARNF_n, FLTOUT, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74LVC06 U13053(STRT2, MOSCAL_n, INKL_n, MINKL, net_U13038_Pad13, MREQIN, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6
endmodule