`timescale 1ns/1ps

module crosspoint_nqi(VCC, GND, SIM_RST, GOJAM, T01, T01_n, T02_n, T03_n, T04_n, T05_n, T06_n, T07_n, T08_n, T09_n, T10_n, T11_n, T12, T12_n, T12USE_n, BR1, BR1_n, BR2, BR2_n, BR12B_n, BR1B2_n, BRDIF_n, S11, S12, INCSET_n, INKL_n, MONPCH, MONWBK, ADS0, CCS0, CCS0_n, CHINC_n, DAS0, DAS0_n, DAS1, DAS1_n, DV1, DV1_n, DV4, DV4_n, DIV_n, DXCH0, FETCH0, FETCH0_n, GOJ1, GOJ1_n, INOUT, INOUT_n, MASK0, MASK0_n, MP0, MP3, MP3_n, MSU0, MSU0_n, NDX0_n, PRINC, QXCH0_n, RAND0, READ0, ROR0, RSM3, RSM3_n, RUPT0, RXOR0, RXOR0_n, SHANC_n, SHIFT, SHIFT_n, STFET1_n, TC0, TC0_n, TCF0, TCSAJ3_n, TS0, TS0_n, WAND0, WOR0, IC1, IC2, IC2_n, IC3, IC4, IC5, IC5_n, IC8_n, IC9, IC10, IC10_n, IC11_n, IC12, IC12_n, IC13, IC14, IC15_n, IC16, IC16_n, C24A, C25A, C26A, C27A, C30A, C37P, C40P, C41P, C42P, C43P, C44P, XT0_n, XT2_n, XT3_n, XT4_n, XT5_n, XT6_n, YB0_n, YT0_n, n5XP9, n5XP11, n10XP6, DVST, NDR100_n, NISQ, RSTSTG, TOV_n, TPZG_n, TRSM);
    input wire SIM_RST;
    input wire ADS0;
    input wire BR1;
    input wire BR12B_n;
    input wire BR1B2_n;
    input wire BR1_n;
    input wire BR2;
    input wire BR2_n;
    input wire BRDIF_n;
    input wire C24A;
    input wire C25A;
    input wire C26A;
    input wire C27A;
    input wire C30A;
    input wire C37P;
    input wire C40P;
    input wire C41P;
    input wire C42P;
    input wire C43P;
    input wire C44P;
    input wire CCS0;
    input wire CCS0_n;
    input wire CHINC_n;
    input wire DAS0;
    input wire DAS0_n;
    input wire DAS1;
    input wire DAS1_n;
    input wire DIV_n;
    input wire DV1;
    input wire DV1_n;
    input wire DV4;
    input wire DV4_n;
    output wire DVST;
    input wire DXCH0;
    input wire FETCH0;
    input wire FETCH0_n;
    input wire GND;
    input wire GOJ1;
    input wire GOJ1_n;
    input wire GOJAM;
    input wire IC1;
    input wire IC10;
    input wire IC10_n;
    input wire IC11_n;
    input wire IC12;
    input wire IC12_n;
    input wire IC13;
    input wire IC14;
    input wire IC15_n;
    input wire IC16;
    input wire IC16_n;
    input wire IC2;
    input wire IC2_n;
    input wire IC3;
    input wire IC4;
    input wire IC5;
    input wire IC5_n;
    input wire IC8_n;
    input wire IC9;
    input wire INCSET_n;
    input wire INKL_n;
    input wire INOUT;
    input wire INOUT_n;
    input wire MASK0;
    input wire MASK0_n;
    input wire MONPCH;
    input wire MONWBK;
    input wire MP0;
    input wire MP3;
    input wire MP3_n;
    input wire MSU0;
    input wire MSU0_n;
    output wire NDR100_n;
    input wire NDX0_n;
    wire NET_206;
    wire NET_207;
    wire NET_208;
    wire NET_209;
    wire NET_210;
    wire NET_211;
    wire NET_212;
    wire NET_213;
    wire NET_214;
    wire NET_215;
    wire NET_216;
    wire NET_217;
    wire NET_220;
    wire NET_222;
    wire NET_223;
    wire NET_224;
    wire NET_225;
    wire NET_227;
    wire NET_228;
    wire NET_229;
    wire NET_230;
    wire NET_231;
    wire NET_232;
    wire NET_233;
    wire NET_236;
    wire NET_237;
    wire NET_238;
    wire NET_239;
    wire NET_240;
    wire NET_241;
    wire NET_242;
    wire NET_243;
    wire NET_244;
    wire NET_245;
    wire NET_246;
    wire NET_247;
    wire NET_248;
    wire NET_249;
    wire NET_250;
    wire NET_251;
    wire NET_252;
    wire NET_253;
    wire NET_254;
    wire NET_255;
    wire NET_256;
    wire NET_257;
    wire NET_258;
    wire NET_259;
    wire NET_260;
    wire NET_261;
    wire NET_262;
    wire NET_263;
    wire NET_264;
    wire NET_265;
    wire NET_266;
    wire NET_267;
    wire NET_269;
    wire NET_270;
    wire NET_271;
    wire NET_272;
    wire NET_273;
    wire NET_274;
    wire NET_275;
    wire NET_276;
    wire NET_277;
    wire NET_278;
    wire NET_279;
    wire NET_280;
    wire NET_281;
    wire NET_282;
    wire NET_283;
    wire NET_284;
    wire NET_285;
    wire NET_287;
    wire NET_288;
    wire NET_289;
    wire NET_290;
    wire NET_291;
    wire NET_292;
    wire NET_293;
    wire NET_294;
    wire NET_295;
    wire NET_296;
    wire NET_297;
    wire NET_298;
    wire NET_299;
    wire NET_300;
    wire NET_301;
    wire NET_302;
    wire NET_303;
    wire NET_304;
    wire NET_305;
    wire NET_306;
    wire NET_307;
    wire NET_308;
    wire NET_310;
    wire NET_311;
    wire NET_312;
    wire NET_313;
    wire NET_314;
    wire NET_315;
    wire NET_316;
    wire NET_317;
    wire NET_318;
    wire NET_320;
    wire NET_322;
    wire NET_324;
    wire NET_325;
    wire NET_326;
    wire NET_327;
    wire NET_328;
    wire NET_329;
    wire NET_330;
    wire NET_331;
    wire NET_333;
    wire NET_335;
    wire NET_336;
    wire NET_337;
    wire NET_338;
    wire NET_339;
    wire NET_340;
    wire NET_341;
    wire NET_342;
    wire NET_344;
    wire NET_345;
    wire NET_347;
    wire NET_348;
    wire NET_349;
    wire NET_350;
    wire NET_351;
    wire NET_352;
    wire NET_353;
    wire NET_354;
    wire NET_355;
    wire NET_358;
    wire NET_359;
    wire NET_361;
    wire NET_362;
    wire NET_363;
    wire NET_364;
    wire NET_365;
    wire NET_366;
    wire NET_367;
    wire NET_368;
    wire NET_369;
    wire NET_370;
    wire NET_371;
    wire NET_372;
    wire NET_373;
    wire NET_374;
    wire NET_375;
    wire NET_376;
    wire NET_377;
    wire NET_378;
    wire NET_379;
    wire NET_380;
    wire NET_381;
    wire NET_382;
    wire NET_383;
    wire NET_384;
    wire NET_385;
    wire NET_386;
    wire NET_387;
    wire NET_388;
    wire NET_389;
    wire NET_390;
    wire NET_391;
    wire NET_392;
    output wire NISQ;
    input wire PRINC;
    input wire QXCH0_n;
    input wire RAND0;
    input wire READ0;
    input wire ROR0;
    input wire RSM3;
    input wire RSM3_n;
    output wire RSTSTG;
    input wire RUPT0;
    input wire RXOR0;
    input wire RXOR0_n;
    input wire S11;
    input wire S12;
    input wire SHANC_n;
    input wire SHIFT;
    input wire SHIFT_n;
    wire STD2;
    input wire STFET1_n;
    input wire T01;
    input wire T01_n;
    input wire T02_n;
    input wire T03_n;
    input wire T04_n;
    input wire T05_n;
    input wire T06_n;
    input wire T07_n;
    input wire T08_n;
    input wire T09_n;
    input wire T10_n;
    input wire T11_n;
    input wire T12;
    input wire T12USE_n;
    input wire T12_n;
    input wire TC0;
    input wire TC0_n;
    input wire TCF0;
    input wire TCSAJ3_n;
    inout wire TOV_n;
    output wire TPZG_n;
    output wire TRSM;
    input wire TS0;
    input wire TS0_n;
    input wire VCC;
    input wire WAND0;
    input wire WOR0;
    input wire XT0_n;
    input wire XT2_n;
    input wire XT3_n;
    input wire XT4_n;
    input wire XT5_n;
    input wire XT6_n;
    input wire YB0_n;
    input wire YT0_n;
    wire __A05_1__10XP1;
    wire __A05_1__10XP7;
    wire __A05_1__10XP8;
    wire __A05_1__11XP2;
    wire __A05_1__2XP7;
    wire __A05_1__3XP5;
    wire __A05_1__3XP6;
    wire __A05_1__4XP5;
    wire __A05_1__5XP12;
    wire __A05_1__7XP4;
    wire __A05_1__7XP9;
    wire __A05_1__8XP12;
    wire __A05_1__8XP15;
    wire __A05_1__8XP3;
    wire __A05_1__9XP5;
    wire __A05_1__A2X_n;
    wire __A05_1__CI_n;
    wire __A05_1__DV1B1B;
    wire __A05_1__GHNHC;
    wire __A05_1__MNISQ;
    wire __A05_1__MONEX_n;
    wire __A05_1__NISQ_n;
    wire __A05_1__PARTC;
    wire __A05_1__PINC;
    wire __A05_1__PINC_n;
    wire __A05_1__PTWOX;
    wire __A05_1__RAD;
    wire __A05_1__RA_n;
    wire __A05_1__RB_n;
    wire __A05_1__RC_n;
    wire __A05_1__RG_n;
    wire __A05_1__RL_n;
    wire __A05_1__RSTRT;
    wire __A05_1__RU_n;
    wire __A05_1__RZ_n;
    wire __A05_1__ST2_n;
    wire __A05_1__TMZ_n;
    wire __A05_1__TSGN_n;
    wire __A05_1__TSUDO_n;
    wire __A05_1__WA_n;
    wire __A05_1__WB_n;
    wire __A05_1__WG_n;
    wire __A05_1__WY12_n;
    wire __A05_1__WY_n;
    wire __A05_1__WZ_n;
    wire __A05_2__10XP10;
    wire __A05_2__11XP6;
    wire __A05_2__2XP8;
    wire __A05_2__5XP13;
    wire __A05_2__5XP15;
    wire __A05_2__5XP19;
    wire __A05_2__5XP21;
    wire __A05_2__6XP2;
    wire __A05_2__6XP7;
    wire __A05_2__6XP8;
    wire __A05_2__A2X_n;
    wire __A05_2__CI_n;
    wire __A05_2__DV4B1B;
    wire __A05_2__OCTAD2;
    wire __A05_2__OCTAD3;
    wire __A05_2__OCTAD4;
    wire __A05_2__OCTAD5;
    wire __A05_2__OCTAD6;
    wire __A05_2__R6;
    wire __A05_2__RA_n;
    wire __A05_2__RB_n;
    wire __A05_2__RC_n;
    wire __A05_2__RG_n;
    wire __A05_2__RL_n;
    wire __A05_2__RQ_n;
    wire __A05_2__RSCT;
    wire __A05_2__RU_n;
    wire __A05_2__RZ_n;
    wire __A05_2__SCAD;
    wire __A05_2__SCAD_n;
    wire __A05_2__TMZ_n;
    wire __A05_2__TSGN_n;
    wire __A05_2__U2BBK;
    wire __A05_2__WA_n;
    wire __A05_2__WB_n;
    wire __A05_2__WL_n;
    wire __A05_2__WS_n;
    wire __A05_2__WY12_n;
    wire __A05_2__WYD_n;
    wire __A05_2__WY_n;
    wire __A05_2__WZ_n;
    wire __A05_2__Z15_n;
    wire __A05_2__Z16_n;
    output wire n10XP6;
    input wire n5XP11;
    output wire n5XP9;

    pullup R5001(NET_227);
    pullup R5002(NET_327);
    pullup R5003(NET_328);
    pullup R5004(__A05_2__RL_n);
    pullup R5005(__A05_2__RA_n);
    pullup R5006(__A05_2__WY_n);
    pullup R5007(__A05_2__WY12_n);
    pullup R5008(__A05_2__SCAD);
    pullup R5009(NET_344);
    pullup R5010(NET_350);
    pullup R5011(__A05_2__TMZ_n);
    U74HC27 U5001(IC10, IC3, TC0, TCF0, IC4, NET_259, GND, NET_258, IC2, IC3, RSM3, NET_261, IC2, VCC, SIM_RST);
    U74HC02 U5002(NET_260, STD2, IC2, NET_282, T01_n, NET_261, GND, T01_n, NET_260, NET_263, IC10_n, T01_n, NET_264, VCC, SIM_RST);
    U74HC02 U5003(NET_279, T01_n, NET_259, NET_262, T02_n, NET_258, GND, T08_n, CCS0_n, NET_211, T02_n, MP3_n, __A05_1__2XP7, VCC, SIM_RST);
    U74HC27 U5004(T02_n, STD2, n10XP6, __A05_1__10XP7, NET_264, NET_267, GND, NET_271, NET_263, __A05_1__3XP6, NET_254, DVST, DIV_n, VCC, SIM_RST);
    U74LVC07 U5005(NET_267, __A05_1__MONEX_n, NET_271, __A05_1__RZ_n, NET_272, __A05_1__RB_n, GND, __A05_1__RA_n, NET_269, __A05_1__WA_n, NET_257, __A05_1__RL_n, NET_251, VCC, SIM_RST);
    U74HC27 U5006(NET_262, __A05_1__8XP15, NET_252, NET_255, __A05_1__8XP12, NET_251, GND, __A05_1__PARTC, INKL_n, SHIFT, MONPCH, __A05_1__NISQ_n, __A05_1__2XP7, VCC, SIM_RST);
    U74HC02 U5007(__A05_1__3XP5, T03_n, IC2_n, NET_288, T01_n, IC15_n, GND, NET_288, NET_270, NET_269, T03_n, TC0_n, __A05_1__3XP6, VCC, SIM_RST);
    U74HC02 U5008(NET_270, T04_n, IC2_n, NET_256, T02_n, IC15_n, GND, NET_256, NET_287, TPZG_n, T04_n, DAS0_n, NET_252, VCC, SIM_RST);
    U74HC02 U5009(NET_257, NET_252, NET_253, NET_253, T04_n, MASK0_n, GND, MP3_n, T10_n, NET_255, T05_n, IC2_n, NET_254, VCC, SIM_RST);
    U74HC02 U5010(NET_287, T05_n, NET_266, NET_265, NET_288, NET_287, GND, T05_n, DAS0_n, __A05_1__5XP12, T06_n, RSM3_n, NET_292, VCC, SIM_RST);
    U74HC27 U5011(__A05_1__PARTC, PRINC, NET_287, NET_288, __A05_1__7XP9, __A05_1__TSGN_n, GND, NET_293, __A05_1__9XP5, NET_288, NET_292, NET_266, CCS0, VCC, SIM_RST);
    U74LVC07 U5012(NET_265, __A05_1__TMZ_n, NET_293, __A05_1__WG_n, NET_290, __A05_1__RG_n, GND, __A05_1__RC_n, NET_291, __A05_1__A2X_n, NET_274, __A05_1__WY_n, NET_276, VCC, SIM_RST);
    U74HC02 U5013(NET_275, T06_n, DAS0_n, NET_289, T06_n, MSU0_n, GND, NET_253, NET_289, NET_291, T07_n, DAS0_n, NET_278, VCC, SIM_RST);
    U74HC27 U5014(NET_287, NET_273, NET_273, NET_275, NET_289, NET_274, GND, NET_276, NET_273, NET_289, NET_275, NET_290, NET_275, VCC, SIM_RST);
    U74HC4002 U5015(NET_272, NET_279, __A05_1__3XP5, NET_278, NET_292, NET_277, GND, NET_280, IC3, RSM3, MP3, IC16, __A05_1__TSUDO_n, VCC, SIM_RST);
    U74HC02 U5016(__A05_1__7XP9, T07_n, MSU0_n, NET_273, T07_n, IC2_n, GND, T07_n, CCS0_n, NET_285, NET_216, NET_206, NET_215, VCC, SIM_RST);
    U74HC27 U5017(NET_289, NET_282, __A05_1__8XP3, NET_285, __A05_1__4XP5, NET_283, GND, NET_281, __A05_1__4XP5, NET_285, NET_282, NET_284, n10XP6, VCC, SIM_RST);
    U74LVC07 U5018(NET_284, __A05_1__CI_n, NET_283, __A05_1__RZ_n, NET_281, __A05_1__WY12_n, GND, __A05_1__WZ_n, NET_217, __A05_1__RB_n, NET_215, __A05_1__WB_n, NET_224, VCC, SIM_RST);
    U74HC27 U5019(CCS0_n, T07_n, BR1_n, CCS0_n, T07_n, __A05_1__PTWOX, GND, NET_217, __A05_1__3XP5, NET_208, NET_211, __A05_1__7XP4, BR2_n, VCC, SIM_RST);
    U74HC27 U5020(INKL_n, FETCH0, NET_211, NET_222, __A05_1__9XP5, NET_210, GND, NET_223, IC2, IC4, DXCH0, NET_216, T08_n, VCC, SIM_RST);
    U74HC02 U5021(__A05_1__RAD, __A05_1__TSUDO_n, T08_n, NET_224, __A05_1__RAD, NET_212, GND, T08_n, NET_225, __A05_1__8XP15, T08_n, NET_220, __A05_1__8XP3, VCC, SIM_RST);
    U74HC04 U5022(IC16, NET_225, NET_301, __A05_2__RQ_n, MP3, NET_312, GND, __A05_2__SCAD_n, __A05_2__SCAD, NDR100_n, NET_306, NET_354, NET_355, VCC, SIM_RST);
    U74HC02 U5023(NET_220, MP0, IC1, NET_222, T08_n, NET_223, GND, T08_n, NET_209, NET_212, T08_n, GOJ1_n, __A05_1__RSTRT, VCC, SIM_RST);
    U74LVC07 U5024(NET_210, __A05_1__RU_n, NET_214, __A05_1__RA_n, NET_213, __A05_1__ST2_n, GND, __A05_1__WY_n, NET_244, __A05_1__RC_n, NET_248, __A05_1__RC_n, NET_232, VCC, SIM_RST);
    U74HC27 U5025(DXCH0, GOJ1, T08_n, BR2, T10_n, n10XP6, GND, NET_245, IC1, IC10, RUPT0, NET_209, DAS0, VCC, SIM_RST);
    U74HC02 U5026(__A05_1__8XP12, T08_n, DAS0_n, NET_208, T08_n, TCSAJ3_n, GND, T09_n, NET_207, NET_206, IC2, __A05_1__DV1B1B, NET_207, VCC, SIM_RST);
    U74HC02 U5027(__A05_1__9XP5, T09_n, DAS0_n, NET_241, T09_n, MASK0_n, GND, NET_241, NET_243, NET_214, T10_n, T08_n, NET_240, VCC, SIM_RST);
    U74HC02 U5028(NET_213, NET_208, NET_240, __A05_1__10XP1, NET_245, T10_n, GND, T10_n, NET_242, NET_243, DAS0, NET_250, NET_242, VCC, SIM_RST);
    U74HC27 U5029(NET_240, NET_241, T10_n, DAS0_n, BR1B2_n, __A05_1__10XP8, GND, NET_232, NET_206, NET_231, n5XP11, NET_244, NET_243, VCC, SIM_RST);
    U74HC02 U5030(NET_250, MSU0_n, BR1_n, __A05_1__10XP7, T10_n, NET_246, GND, NET_250, NET_249, NET_246, BR12B_n, DAS0_n, NET_249, VCC, SIM_RST);
    U74HC02 U5031(__A05_1__11XP2, T11_n, MSU0_n, NET_247, T10_n, MASK0_n, GND, NET_241, NET_247, NET_248, T10_n, NET_233, NET_231, VCC, SIM_RST);
    U74HC02 U5032(NET_233, MSU0, IC14, NET_238, INCSET_n, NET_227, GND, GOJAM, __A05_1__GHNHC, NET_239, NET_239, T01, __A05_1__GHNHC, VCC, SIM_RST);
    U74HC4002 U5033(NET_229, C24A, C25A, C26A, C27A, NET_237, GND, NET_236, C30A, C37P, C40P, C41P, NET_228, VCC, SIM_RST);
    U74HC27 U5034(C42P, C43P, IC12, DAS0, DAS1, NET_374, GND, NET_370, NET_326, NET_325, __A05_2__RSCT, NET_230, C44P, VCC, SIM_RST);
    U74LVC07 U5035(NET_229, NET_227, NET_228, NET_227, NET_230, NET_227, GND, NET_327, NET_374, NET_327, NET_373, __A05_2__WS_n, NET_370, VCC, SIM_RST);
    U74HC02 U5036(__A05_1__PINC_n, NET_238, __A05_1__PINC, __A05_1__PINC, __A05_1__PINC_n, T12, GND, T01_n, NET_327, NET_326, T01_n, FETCH0_n, __A05_2__R6, VCC, SIM_RST);
    U74HC4002 U5037(NET_373, IC9, DXCH0, PRINC, INOUT, NET_372, GND, NET_371, YB0_n, YT0_n, S12, S11, NET_306, VCC, SIM_RST);
    U74HC02 U5038(NET_325, T01_n, CHINC_n, NET_304, T03_n, NET_328, GND, IC5, MP0, NET_375, T03_n, IC8_n, NET_302, VCC, SIM_RST);
    U74HC27 U5039(T01_n, MONPCH, TS0, DAS0, MASK0, NET_378, GND, NET_376, NET_304, NET_302, NET_301, __A05_2__RSCT, INKL_n, VCC, SIM_RST);
    wire U5040_3_NC;
    wire U5040_4_NC;
    wire U5040_5_NC;
    wire U5040_6_NC;
    wire U5040_8_NC;
    wire U5040_9_NC;
    wire U5040_10_NC;
    wire U5040_11_NC;
    U74HC27 U5040(NET_305, NET_296, U5040_3_NC, U5040_4_NC, U5040_5_NC, U5040_6_NC, GND, U5040_8_NC, U5040_9_NC, U5040_10_NC, U5040_11_NC, NET_377, __A05_2__6XP2, VCC, SIM_RST);
    U74LVC07 U5041(NET_376, __A05_2__WB_n, NET_377, __A05_2__WB_n, NET_378, NET_328, GND, NET_328, NET_375, __A05_2__RL_n, NET_365, __A05_2__RA_n, NET_366, VCC, SIM_RST);
    U74HC02 U5042(__A05_2__2XP8, T02_n, FETCH0_n, NET_301, T03_n, QXCH0_n, GND, T04_n, DV1_n, NET_300, T04_n, NET_303, NET_305, VCC, SIM_RST);
    U74HC27 U5043(NET_302, NET_300, DV1, INOUT, IC2, NET_303, GND, NET_364, NET_296, NET_295, n5XP9, NET_365, __A05_2__11XP6, VCC, SIM_RST);
    U74HC02 U5044(NET_366, NET_304, __A05_2__6XP2, TRSM, T05_n, NDX0_n, GND, IC12_n, NET_294, NET_296, DAS1_n, NET_310, NET_295, VCC, SIM_RST);
    U74HC27 U5045(__A05_2__5XP13, __A05_2__5XP15, DAS1, PRINC, __A05_1__PARTC, NET_298, GND, NET_369, NET_299, __A05_2__2XP8, __A05_2__10XP10, NET_363, NET_307, VCC, SIM_RST);
    U74LVC07 U5046(NET_364, __A05_2__RG_n, NET_363, __A05_2__RG_n, NET_369, __A05_2__WY_n, GND, __A05_2__A2X_n, NET_367, __A05_2__CI_n, NET_368, __A05_2__WY12_n, NET_389, VCC, SIM_RST);
    U74HC02 U5047(NET_299, NET_298, NET_310, NET_367, NET_295, __A05_2__10XP10, GND, SHIFT_n, NET_310, n5XP9, SHANC_n, NET_310, NET_297, VCC, SIM_RST);
    U74HC27 U5048(NET_297, NET_313, YT0_n, YB0_n, XT0_n, NET_392, GND, NET_349, RAND0, WAND0, NET_355, NET_368, NET_311, VCC, SIM_RST);
    U74HC02 U5049(__A05_2__5XP13, IC8_n, NET_310, __A05_2__5XP15, QXCH0_n, NET_310, GND, NET_308, NET_310, __A05_2__5XP21, IC5_n, NET_310, NET_307, VCC, SIM_RST);
    U74HC02 U5050(NET_313, IC16_n, NET_310, NET_311, NET_312, NET_310, GND, NET_313, NET_311, NET_389, S11, S12, NET_390, VCC, SIM_RST);
    U74LVC07 U5051(NET_388, __A05_2__RB_n, NET_391, __A05_2__RZ_n, NET_390, __A05_2__SCAD, GND, __A05_2__SCAD, NET_392, __A05_2__RC_n, NET_381, NET_344, NET_379, VCC, SIM_RST);
    U74HC02 U5052(NET_388, __A05_2__5XP19, NET_313, NET_391, __A05_2__6XP7, NET_311, GND, XT2_n, NDR100_n, __A05_2__OCTAD2, NDR100_n, XT3_n, __A05_2__OCTAD3, VCC, SIM_RST);
    U74HC02 U5053(__A05_2__OCTAD4, NDR100_n, XT4_n, __A05_2__OCTAD5, NDR100_n, XT5_n, GND, NDR100_n, XT6_n, __A05_2__OCTAD6, BR1_n, DV1_n, NET_355, VCC, SIM_RST);
    U74HC02 U5054(NET_348, NET_349, T05_n, __A05_2__5XP19, T05_n, NET_347, GND, DV1_n, BR1, __A05_1__DV1B1B, TS0_n, BRDIF_n, NET_345, VCC, SIM_RST);
    U74HC4002 U5055(NET_381, NET_348, NET_351, NET_341, NET_342, NET_383, GND, NET_382, __A05_2__5XP13, NET_316, NET_359, NET_336, NET_361, VCC, SIM_RST);
    U74HC27 U5056(ROR0, __A05_1__DV1B1B, IC2, IC5, READ0, NET_379, GND, NET_384, IC2, IC3, TS0, NET_347, WOR0, VCC, SIM_RST);
    U74HC02 U5057(NET_380, NET_345, DV4, NET_352, NET_344, T05_n, GND, NET_354, T05_n, NET_353, NET_352, NET_351, NET_386, VCC, SIM_RST);
    U74LVC07 U5058(NET_380, NET_344, NET_387, __A05_2__Z16_n, NET_386, __A05_2__WA_n, GND, NET_350, NET_384, NET_350, NET_385, __A05_2__WZ_n, NET_322, VCC, SIM_RST);
    U74HC04 U5059(NET_353, NET_387, NET_324, NET_322, NET_351, NET_358, GND, NET_339, NET_341, NISQ, __A05_1__NISQ_n, __A05_1__MNISQ, __A05_1__NISQ_n, VCC, SIM_RST);
    U74HC02 U5060(NET_385, IC16, MP3, NET_324, T06_n, NET_350, GND, T06_n, DAS1_n, __A05_2__6XP8, __A05_2__6XP8, __A05_2__6XP7, NET_320, VCC, SIM_RST);
    U74LVC07 U5061(NET_320, TOV_n, NET_315, __A05_2__RU_n, NET_314, __A05_2__RU_n, GND, __A05_2__WB_n, NET_331, __A05_2__RG_n, NET_330, __A05_2__TSGN_n, NET_362, VCC, SIM_RST);
    U74HC02 U5062(__A05_2__6XP7, DV4_n, T06_n, NET_329, T07_n, NET_318, GND, T07_n, STFET1_n, NET_333, T08_n, DV4_n, RSTSTG, VCC, SIM_RST);
    U74HC27 U5063(NET_324, __A05_2__6XP8, NET_317, NET_359, NET_316, NET_314, GND, __A05_2__6XP2, T06_n, RXOR0, INOUT_n, NET_315, n5XP11, VCC, SIM_RST);
    U74HC27 U5064(IC13, IC14, NET_329, NET_359, NET_317, NET_331, GND, NET_330, NET_329, NET_333, NET_342, NET_318, DV1, VCC, SIM_RST);
    U74HC27 U5065(T08_n, MONWBK, IC2, IC14, DV1, NET_335, GND, NET_337, __A05_2__DV4B1B, IC4, NET_338, __A05_2__U2BBK, STFET1_n, VCC, SIM_RST);
    U74HC02 U5066(NET_362, RSTSTG, n5XP9, NET_351, T09_n, NET_354, GND, T09_n, DV4_n, NET_359, T09_n, DAS1_n, NET_341, VCC, SIM_RST);
    wire U5067_10_NC;
    wire U5067_11_NC;
    wire U5067_12_NC;
    wire U5067_13_NC;
    U74LVC07 U5067(NET_358, __A05_2__Z15_n, NET_361, __A05_2__WL_n, NET_339, __A05_2__TMZ_n, GND, __A05_2__WYD_n, NET_340, U5067_10_NC, U5067_11_NC, U5067_12_NC, U5067_13_NC, VCC, SIM_RST);
    wire U5068_4_NC;
    wire U5068_5_NC;
    wire U5068_6_NC;
    U74HC02 U5068(NET_317, T10_n, NET_335, U5068_4_NC, U5068_5_NC, U5068_6_NC, GND, T10_n, IC11_n, __A05_2__10XP10, T10_n, NET_337, NET_336, VCC, SIM_RST);
    wire U5069_8_NC;
    wire U5069_9_NC;
    wire U5069_10_NC;
    wire U5069_11_NC;
    U74HC27 U5069(DAS1_n, ADS0, T12_n, T12USE_n, DV1_n, NET_316, GND, U5069_8_NC, U5069_9_NC, U5069_10_NC, U5069_11_NC, NET_338, BR2, VCC, SIM_RST);
    U74HC02 U5070(__A05_2__DV4B1B, DV4_n, BR1, __A05_2__11XP6, T11_n, DV1_n, GND, n5XP9, __A05_2__11XP6, NET_340, T11_n, RXOR0_n, NET_342, VCC, SIM_RST);
endmodule