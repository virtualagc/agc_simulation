`timescale 1ns/1ps

module parity_s_register(VCC, GND, SIM_RST, GOJAM, PHS4_n, T02_n, T07_n, T12A, TPARG_n, TSUDO_n, FUTEXT, CGG, CSG, WEDOPG_n, WSG_n, G01, G02, G03, G04, G05, G06, G07, G08, G09, G10, G11, G12, G13, G14, G15, G16, WL01_n, WL02_n, WL03_n, WL04_n, WL05_n, WL06_n, WL07_n, WL08_n, WL09_n, WL10_n, WL11_n, WL12_n, WL13_n, WL14_n, RAD, SAP, SCAD, OCTAD2, n8XP5, MONPAR, XB0_n, XB1_n, XB2_n, XB3_n, CYL_n, CYR_n, EDOP_n, GINH, SR_n, EXTPLS, INHPLS, RELPLS, G01ED, G02ED, G03ED, G04ED, G05ED, G06ED, G07ED, GEQZRO_n, RADRG, RADRZ, S11, S12);
    input wire SIM_RST;
    input wire CGG;
    input wire CSG;
    output wire CYL_n;
    output wire CYR_n;
    output wire EDOP_n;
    output wire EXTPLS;
    input wire FUTEXT;
    input wire G01;
    output wire G01ED;
    input wire G02;
    output wire G02ED;
    input wire G03;
    output wire G03ED;
    input wire G04;
    output wire G04ED;
    input wire G05;
    output wire G05ED;
    input wire G06;
    output wire G06ED;
    input wire G07;
    output wire G07ED;
    input wire G08;
    input wire G09;
    input wire G10;
    input wire G11;
    input wire G12;
    input wire G13;
    input wire G14;
    input wire G15;
    input wire G16;
    output wire GEQZRO_n;
    output wire GINH;
    input wire GND;
    input wire GOJAM;
    inout wire INHPLS;
    input wire MONPAR;
    wire NET_106;
    wire NET_107;
    wire NET_108;
    wire NET_109;
    wire NET_110;
    wire NET_111;
    wire NET_112;
    wire NET_113;
    wire NET_114;
    wire NET_116;
    wire NET_118;
    wire NET_119;
    wire NET_120;
    wire NET_121;
    wire NET_122;
    wire NET_123;
    wire NET_124;
    wire NET_125;
    wire NET_126;
    wire NET_127;
    wire NET_128;
    wire NET_129;
    wire NET_130;
    wire NET_131;
    wire NET_132;
    wire NET_133;
    wire NET_134;
    wire NET_135;
    wire NET_136;
    wire NET_137;
    wire NET_138;
    wire NET_139;
    wire NET_140;
    wire NET_141;
    wire NET_142;
    wire NET_143;
    wire NET_146;
    wire NET_147;
    wire NET_148;
    wire NET_149;
    wire NET_150;
    wire NET_151;
    wire NET_155;
    wire NET_156;
    wire NET_165;
    wire NET_166;
    wire NET_168;
    wire NET_172;
    wire NET_173;
    wire NET_174;
    wire NET_177;
    wire NET_178;
    wire NET_179;
    wire NET_180;
    wire NET_181;
    wire NET_182;
    wire NET_183;
    wire NET_184;
    wire NET_185;
    wire NET_186;
    wire NET_189;
    wire NET_190;
    wire NET_191;
    wire NET_192;
    wire NET_193;
    wire NET_194;
    wire NET_195;
    wire NET_196;
    wire NET_197;
    wire NET_198;
    wire NET_199;
    wire NET_200;
    wire NET_204;
    wire NET_205;
    wire NET_206;
    wire NET_207;
    wire NET_208;
    wire NET_209;
    wire NET_210;
    wire NET_211;
    wire NET_212;
    wire NET_213;
    wire NET_214;
    wire NET_215;
    wire NET_216;
    wire NET_217;
    wire NET_218;
    wire NET_219;
    wire NET_220;
    wire NET_221;
    wire NET_222;
    wire NET_223;
    wire NET_224;
    wire NET_225;
    wire NET_226;
    wire NET_227;
    wire NET_228;
    wire NET_229;
    wire NET_230;
    wire NET_231;
    wire NET_232;
    wire NET_233;
    wire NET_234;
    wire NET_235;
    wire NET_236;
    wire NET_237;
    wire NET_238;
    wire NET_239;
    wire NET_240;
    wire NET_241;
    wire NET_242;
    wire NET_243;
    wire NET_244;
    wire NET_245;
    wire NET_246;
    wire NET_247;
    wire NET_248;
    wire NET_249;
    wire NET_250;
    wire NET_251;
    wire NET_252;
    input wire OCTAD2;
    input wire PHS4_n;
    input wire RAD;
    output wire RADRG;
    output wire RADRZ;
    inout wire RELPLS;
    output wire S11;
    output wire S12;
    input wire SAP;
    input wire SCAD;
    output wire SR_n;
    input wire T02_n;
    input wire T07_n;
    input wire T12A;
    input wire TPARG_n;
    input wire TSUDO_n;
    input wire VCC;
    input wire WEDOPG_n;
    input wire WL01_n;
    input wire WL02_n;
    input wire WL03_n;
    input wire WL04_n;
    input wire WL05_n;
    input wire WL06_n;
    input wire WL07_n;
    input wire WL08_n;
    input wire WL09_n;
    input wire WL10_n;
    input wire WL11_n;
    input wire WL12_n;
    input wire WL13_n;
    input wire WL14_n;
    input wire WSG_n;
    input wire XB0_n;
    input wire XB1_n;
    input wire XB2_n;
    input wire XB3_n;
    wire __A12_1__G01A_n;
    wire __A12_1__G02_n;
    wire __A12_1__G03_n;
    wire __A12_1__GEMP;
    wire __A12_1__GNZRO;
    wire __A12_1__MGP_n;
    wire __A12_1__MPAL;
    wire __A12_1__MSP;
    wire __A12_1__PA03;
    wire __A12_1__PA03_n;
    wire __A12_1__PA06;
    wire __A12_1__PA06_n;
    wire __A12_1__PA09;
    wire __A12_1__PA09_n;
    wire __A12_1__PA12;
    wire __A12_1__PA12_n;
    wire __A12_1__PA15;
    wire __A12_1__PA15_n;
    wire __A12_1__PALE;
    wire __A12_1__PB09;
    wire __A12_1__PB09_n;
    wire __A12_1__PB15;
    wire __A12_1__PB15_n;
    wire __A12_1__PC15;
    wire __A12_1__PC15_n;
    wire __A12_1__T7PHS4;
    wire __A12_1__T7PHS4_n;
    wire __A12_2__S01;
    wire __A12_2__S01_n;
    wire __A12_2__S02;
    wire __A12_2__S02_n;
    wire __A12_2__S03;
    wire __A12_2__S03_n;
    wire __A12_2__S04;
    wire __A12_2__S04_n;
    wire __A12_2__S05;
    wire __A12_2__S05_n;
    wire __A12_2__S06;
    wire __A12_2__S06_n;
    wire __A12_2__S07;
    wire __A12_2__S07_n;
    wire __A12_2__S08;
    wire __A12_2__S08_n;
    wire __A12_2__S09;
    wire __A12_2__S09_n;
    wire __A12_2__S10;
    wire __A12_2__S10_n;
    wire __A12_2__S11_n;
    wire __A12_2__S12_n;
    input wire n8XP5;

    pullup R12001(__A12_1__GNZRO);
    pullup R12002(RELPLS);
    pullup R12003(INHPLS);
    pullup R12004(__A12_1__PALE);
    U74HC04 U12001(G01, __A12_1__G01A_n, G02, __A12_1__G02_n, G03, __A12_1__G03_n, GND, __A12_1__PA03_n, __A12_1__PA03, NET_196, G04, NET_190, G05, VCC, SIM_RST);
    U74HC27 U12002(G01, G02, G01, __A12_1__G02_n, __A12_1__G03_n, NET_182, GND, NET_181, __A12_1__G01A_n, G02, __A12_1__G03_n, NET_177, G03, VCC, SIM_RST);
    U74HC27 U12003(__A12_1__G01A_n, __A12_1__G02_n, G04, G05, G06, NET_183, GND, NET_186, G04, NET_190, NET_195, NET_180, G03, VCC, SIM_RST);
    U74HC4002 U12004(__A12_1__PA03, NET_177, NET_182, NET_181, NET_180, NET_179, GND, NET_178, NET_183, NET_186, NET_185, NET_184, __A12_1__PA06, VCC, SIM_RST);
    U74HC04 U12005(G06, NET_195, NET_183, NET_133, __A12_1__PA06, __A12_1__PA06_n, GND, NET_189, G07, NET_127, G08, NET_174, G09, VCC, SIM_RST);
    U74HC27 U12006(NET_196, G05, NET_196, NET_190, G06, NET_184, GND, NET_123, G07, G08, G09, NET_185, NET_195, VCC, SIM_RST);
    U74HC27 U12007(G07, NET_127, NET_189, G08, NET_174, NET_126, GND, NET_125, NET_189, NET_127, G09, NET_122, NET_174, VCC, SIM_RST);
    U74HC4002 U12008(__A12_1__PA09, NET_123, NET_122, NET_126, NET_125, NET_173, GND, NET_172, NET_136, NET_135, NET_138, NET_137, __A12_1__PA12, VCC, SIM_RST);
    U74HC04 U12009(NET_123, NET_132, __A12_1__PA09, __A12_1__PA09_n, G10, NET_120, GND, NET_124, G11, NET_121, G12, NET_114, NET_136, VCC, SIM_RST);
    U74HC27 U12010(G10, G11, G10, NET_124, NET_121, NET_135, GND, NET_138, NET_120, G11, NET_121, NET_136, G12, VCC, SIM_RST);
    U74HC27 U12011(NET_120, NET_124, G13, G14, G16, NET_134, GND, NET_130, G13, NET_131, NET_139, NET_137, G12, VCC, SIM_RST);
    U74HC04 U12012(__A12_1__PA12, __A12_1__PA12_n, G13, NET_140, G14, NET_131, GND, NET_139, G16, NET_113, NET_134, __A12_1__PA15_n, __A12_1__PA15, VCC, SIM_RST);
    U74HC27 U12013(NET_140, G14, NET_140, NET_131, G16, NET_128, GND, NET_198, NET_133, NET_132, NET_114, NET_129, NET_139, VCC, SIM_RST);
    U74HC4002 #(0, 1) U12014(__A12_1__PA15, NET_134, NET_130, NET_129, NET_128, NET_200, GND, NET_199, EXTPLS, RELPLS, INHPLS, NET_118, NET_119, VCC, SIM_RST);
    U74HC02 U12015(NET_197, NET_113, G15, NET_110, TSUDO_n, __A12_1__T7PHS4_n, GND, __A12_1__G02_n, G03, NET_192, G02, __A12_1__G03_n, NET_191, VCC, SIM_RST);
    U74LVC07 U12016(NET_198, __A12_1__GNZRO, NET_197, __A12_1__GNZRO, NET_193, RELPLS, GND, RELPLS, NET_192, INHPLS, NET_194, INHPLS, NET_191, VCC, SIM_RST);
    U74HC04 U12017(__A12_1__GNZRO, NET_109, NET_182, NET_112, NET_110, NET_111, GND, GEQZRO_n, NET_108, NET_116, RAD, __A12_1__PB09_n, __A12_1__PB09, VCC, SIM_RST);
    U74HC27 U12018(NET_112, NET_109, NET_109, NET_111, __A12_1__G01A_n, NET_193, GND, NET_194, NET_109, G01, NET_111, EXTPLS, NET_111, VCC, SIM_RST);
    U74HC4002 U12019(NET_108, NET_109, G02, G01, G03, NET_107, GND, NET_106, NET_151, NET_150, NET_149, NET_165, __A12_1__PB09, VCC, SIM_RST);
    U74HC02 U12020(NET_118, NET_119, T12A, RADRZ, NET_119, NET_116, GND, NET_116, NET_118, RADRG, __A12_1__PA12, __A12_1__PA15, NET_156, VCC, SIM_RST);
    U74HC27 U12021(__A12_1__PA03, __A12_1__PA06, __A12_1__PA03, __A12_1__PA06_n, __A12_1__PA09_n, NET_150, GND, NET_149, __A12_1__PA03_n, __A12_1__PA06, __A12_1__PA09_n, NET_151, __A12_1__PA09, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U12022(__A12_1__PA03_n, __A12_1__PA06_n, NET_142, MONPAR, SAP, NET_143, GND, NET_148, SCAD, NET_141, GOJAM, NET_165, __A12_1__PA09, VCC, SIM_RST);
    wire U12023_8_NC;
    wire U12023_9_NC;
    wire U12023_10_NC;
    U74HC02 U12023(NET_155, __A12_1__PA12_n, __A12_1__PA15_n, __A12_1__PB15, NET_156, NET_155, GND, U12023_8_NC, U12023_9_NC, U12023_10_NC, __A12_1__PB09, __A12_1__PB15_n, NET_168, VCC, SIM_RST);
    U74HC04 U12024(__A12_1__PB15, __A12_1__PB15_n, __A12_1__PC15, __A12_1__PC15_n, __A12_1__PC15, __A12_1__MGP_n, GND, __A12_1__GEMP, __A12_1__PC15_n, __A12_1__MSP, NET_143, __A12_1__MPAL, __A12_1__PALE, VCC, SIM_RST);
    U74HC02 U12025(__A12_1__PC15, NET_166, NET_168, NET_142, CGG, NET_143, GND, __A12_1__PC15, NET_142, NET_141, __A12_1__PC15_n, NET_143, NET_146, VCC, SIM_RST);
    U74HC27 U12026(TPARG_n, n8XP5, T07_n, PHS4_n, FUTEXT, __A12_1__T7PHS4, GND, NET_243, XB0_n, T02_n, NET_242, NET_147, NET_146, VCC, SIM_RST);
    wire U12027_5_NC;
    wire U12027_6_NC;
    wire U12027_8_NC;
    wire U12027_9_NC;
    wire U12027_10_NC;
    wire U12027_11_NC;
    wire U12027_12_NC;
    wire U12027_13_NC;
    U74LVC07 U12027(NET_148, __A12_1__PALE, NET_147, __A12_1__PALE, U12027_5_NC, U12027_6_NC, GND, U12027_8_NC, U12027_9_NC, U12027_10_NC, U12027_11_NC, U12027_12_NC, U12027_13_NC, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U12028(G01ED, WEDOPG_n, WL08_n, NET_233, WL08_n, WSG_n, GND, NET_233, NET_232, NET_231, NET_231, CSG, NET_232, VCC, SIM_RST);
    U74HC04 U12029(NET_231, __A12_2__S08, NET_232, __A12_2__S08_n, NET_226, __A12_2__S09, GND, __A12_2__S09_n, NET_225, __A12_2__S10, NET_229, __A12_2__S10_n, NET_228, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U12030(G02ED, WEDOPG_n, WL09_n, NET_227, WL09_n, WSG_n, GND, NET_227, NET_225, NET_226, NET_226, CSG, NET_225, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U12031(G03ED, WEDOPG_n, WL10_n, NET_230, WL10_n, WSG_n, GND, NET_230, NET_228, NET_229, NET_229, CSG, NET_228, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U12032(G04ED, WEDOPG_n, WL11_n, NET_239, WL11_n, WSG_n, GND, NET_239, NET_237, NET_238, NET_238, CSG, NET_237, VCC, SIM_RST);
    U74HC04 U12033(NET_238, S11, NET_237, __A12_2__S11_n, NET_235, S12, GND, __A12_2__S12_n, NET_236, __A12_2__S01, NET_213, __A12_2__S01_n, NET_211, VCC, SIM_RST);
    U74HC02 U12034(G05ED, WEDOPG_n, WL12_n, NET_234, WL12_n, WSG_n, GND, EDOP_n, T12A, NET_250, NET_235, CSG, NET_236, VCC, SIM_RST);
    U74HC02 #(0, 0, 0, 1) U12035(G06ED, WEDOPG_n, WL13_n, G07ED, WEDOPG_n, WL14_n, GND, WL01_n, WSG_n, NET_212, NET_212, NET_211, NET_213, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U12036(NET_211, NET_213, CSG, NET_206, WL02_n, WSG_n, GND, NET_206, NET_205, NET_204, NET_204, CSG, NET_205, VCC, SIM_RST);
    U74HC04 U12037(NET_204, __A12_2__S02, NET_205, __A12_2__S02_n, NET_209, __A12_2__S03, GND, __A12_2__S03_n, NET_208, __A12_2__S04, NET_220, __A12_2__S04_n, NET_222, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U12038(NET_207, WL03_n, WSG_n, NET_209, NET_207, NET_208, GND, NET_209, CSG, NET_208, WL04_n, WSG_n, NET_210, VCC, SIM_RST);
    U74HC02 #(1, 0, 0, 1) U12039(NET_220, NET_210, NET_222, NET_222, NET_220, CSG, GND, WL05_n, WSG_n, NET_223, NET_223, NET_219, NET_221, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U12040(NET_219, NET_221, CSG, NET_224, WL06_n, WSG_n, GND, NET_224, NET_217, NET_218, NET_218, NET_252, NET_217, VCC, SIM_RST);
    U74HC04 U12041(NET_221, __A12_2__S05, NET_219, __A12_2__S05_n, NET_218, __A12_2__S06, GND, __A12_2__S06_n, NET_217, __A12_2__S07, NET_216, __A12_2__S07_n, NET_214, VCC, SIM_RST);
    wire U12042_11_NC;
    wire U12042_12_NC;
    wire U12042_13_NC;
    U74HC02 #(0, 1, 0, 0) U12042(NET_215, WL07_n, WSG_n, NET_216, NET_215, NET_214, GND, NET_216, CSG, NET_214, U12042_11_NC, U12042_12_NC, U12042_13_NC, VCC, SIM_RST);
    wire U12043_3_NC;
    wire U12043_4_NC;
    wire U12043_10_NC;
    wire U12043_11_NC;
    wire U12043_12_NC;
    wire U12043_13_NC;
    U74HC04 U12043(__A12_1__T7PHS4, __A12_1__T7PHS4_n, U12043_3_NC, U12043_4_NC, OCTAD2, NET_242, GND, GINH, NET_249, U12043_10_NC, U12043_11_NC, U12043_12_NC, U12043_13_NC, VCC, SIM_RST);
    wire U12044_1_NC;
    wire U12044_2_NC;
    wire U12044_3_NC;
    wire U12044_4_NC;
    wire U12044_5_NC;
    U74HC4002 U12044(U12044_1_NC, U12044_2_NC, U12044_3_NC, U12044_4_NC, U12044_5_NC, NET_247, GND, NET_248, NET_244, NET_246, NET_245, NET_250, NET_249, VCC, SIM_RST);
    wire U12046_1_NC;
    wire U12046_2_NC;
    wire U12046_3_NC;
    U74HC02 #(0, 1, 0, 1) U12046(U12046_1_NC, U12046_2_NC, U12046_3_NC, CYR_n, NET_243, NET_244, GND, CYR_n, T12A, NET_244, NET_240, NET_246, SR_n, VCC, SIM_RST);
    U74HC27 U12047(NET_242, T02_n, NET_242, T02_n, XB2_n, NET_241, GND, NET_251, NET_242, T02_n, XB3_n, NET_240, XB1_n, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 1) U12048(NET_246, SR_n, T12A, CYL_n, NET_241, NET_245, GND, CYL_n, T12A, NET_245, NET_251, NET_250, EDOP_n, VCC, SIM_RST);
    wire U12049_3_NC;
    wire U12049_4_NC;
    wire U12049_5_NC;
    wire U12049_6_NC;
    wire U12049_8_NC;
    wire U12049_9_NC;
    wire U12049_10_NC;
    wire U12049_11_NC;
    U74HC27 #(1, 0, 0) U12049(n8XP5, NET_234, U12049_3_NC, U12049_4_NC, U12049_5_NC, U12049_6_NC, GND, U12049_8_NC, U12049_9_NC, U12049_10_NC, U12049_11_NC, NET_235, NET_236, VCC, SIM_RST);
    wire U2023_1_NC;
    wire U2023_2_NC;
    wire U2023_3_NC;
    wire U2023_4_NC;
    wire U2023_5_NC;
    wire U2023_6_NC;
    wire U2023_11_NC;
    wire U2023_12_NC;
    wire U2023_13_NC;
    U74HC02 U2023(U2023_1_NC, U2023_2_NC, U2023_3_NC, U2023_4_NC, U2023_5_NC, U2023_6_NC, GND, __A12_1__PB09_n, __A12_1__PB15, NET_166, U2023_11_NC, U2023_12_NC, U2023_13_NC, VCC, SIM_RST);
endmodule