`timescale 1ns/1ps

module four_bit_4(VCC, GND, SIM_RST, A2XG_n, CAG, CBG, CGG, CLG1G, CLXC, CQG, CUG, CZG, L2GDG_n, RAG_n, RCG_n, RGG_n, RLG_n, RQG_n, RZG_n, WAG_n, WALSG_n, WBG_n, WLG_n, WQG_n, WZG_n, CI13_n, CO14, BXVX, MONEX, XUY01_n, XUY02_n, CH13, CH14, CH16, L12_n, G2LSG_n, WL01_n, WL02_n, G01_n, MDT13, MDT14, MDT15, MDT16, SA13, SA14, SA16, RBHG_n, RULOG_n, RUG_n, G16SW_n, WG1G_n, WG2G_n, WG3G_n, WG4G_n, WG5G_n, WYDG_n, WYHIG_n, R1C, US2SG, WL12_n, WHOMPA, EAC_n, G13_n, G14_n, G15_n, L15_n, SUMA15_n, SUMB15_n, SUMA16_n, SUMB16_n, WL13_n, WL14_n, WL15, WL15_n, WL16, WL16_n, XUY13_n, XUY14_n);
    input wire SIM_RST;
    input wire A2XG_n;
    input wire BXVX;
    input wire CAG;
    input wire CBG;
    input wire CGG;
    input wire CH13;
    input wire CH14;
    input wire CH16;
    input wire CI13_n;
    input wire CLG1G;
    input wire CLXC;
    input wire CO14;
    input wire CQG;
    input wire CUG;
    input wire CZG;
    output wire EAC_n;
    input wire G01_n;
    inout wire G13_n;
    inout wire G14_n;
    inout wire G15_n;
    input wire G16SW_n;
    input wire G2LSG_n;
    input wire GND;
    input wire L12_n;
    inout wire L15_n;
    input wire L2GDG_n;
    input wire MDT13;
    input wire MDT14;
    input wire MDT15;
    input wire MDT16;
    input wire MONEX;
    wire NET_129;
    wire NET_130;
    wire NET_131;
    wire NET_132;
    wire NET_133;
    wire NET_134;
    wire NET_135;
    wire NET_136;
    wire NET_137;
    wire NET_138;
    wire NET_139;
    wire NET_140;
    wire NET_141;
    wire NET_144;
    wire NET_147;
    wire NET_148;
    wire NET_149;
    wire NET_150;
    wire NET_151;
    wire NET_152;
    wire NET_153;
    wire NET_154;
    wire NET_155;
    wire NET_156;
    wire NET_159;
    wire NET_160;
    wire NET_161;
    wire NET_162;
    wire NET_165;
    wire NET_166;
    wire NET_167;
    wire NET_168;
    wire NET_169;
    wire NET_170;
    wire NET_171;
    wire NET_172;
    wire NET_173;
    wire NET_174;
    wire NET_175;
    wire NET_176;
    wire NET_177;
    wire NET_178;
    wire NET_179;
    wire NET_180;
    wire NET_181;
    wire NET_182;
    wire NET_183;
    wire NET_184;
    wire NET_185;
    wire NET_186;
    wire NET_187;
    wire NET_188;
    wire NET_189;
    wire NET_190;
    wire NET_191;
    wire NET_192;
    wire NET_197;
    wire NET_198;
    wire NET_199;
    wire NET_201;
    wire NET_202;
    wire NET_203;
    wire NET_204;
    wire NET_205;
    wire NET_206;
    wire NET_207;
    wire NET_208;
    wire NET_209;
    wire NET_210;
    wire NET_211;
    wire NET_212;
    wire NET_213;
    wire NET_214;
    wire NET_215;
    wire NET_216;
    wire NET_217;
    wire NET_218;
    wire NET_219;
    wire NET_220;
    wire NET_221;
    wire NET_222;
    wire NET_223;
    wire NET_224;
    wire NET_225;
    wire NET_226;
    wire NET_227;
    wire NET_228;
    wire NET_229;
    wire NET_230;
    wire NET_231;
    wire NET_232;
    wire NET_233;
    wire NET_234;
    wire NET_237;
    wire NET_240;
    wire NET_241;
    wire NET_242;
    wire NET_243;
    wire NET_244;
    wire NET_245;
    wire NET_246;
    wire NET_247;
    wire NET_248;
    wire NET_249;
    wire NET_252;
    wire NET_253;
    wire NET_254;
    wire NET_255;
    wire NET_258;
    wire NET_259;
    wire NET_260;
    wire NET_261;
    wire NET_262;
    wire NET_263;
    wire NET_264;
    wire NET_265;
    wire NET_266;
    wire NET_267;
    wire NET_268;
    wire NET_269;
    wire NET_270;
    wire NET_271;
    wire NET_272;
    wire NET_273;
    wire NET_274;
    wire NET_275;
    wire NET_276;
    wire NET_277;
    wire NET_278;
    wire NET_279;
    wire NET_280;
    wire NET_281;
    wire NET_282;
    wire NET_283;
    wire NET_285;
    wire NET_286;
    wire NET_290;
    wire NET_291;
    wire NET_292;
    wire NET_294;
    wire NET_295;
    wire NET_296;
    wire NET_297;
    wire NET_298;
    wire NET_299;
    wire NET_300;
    wire NET_301;
    wire NET_302;
    wire NET_303;
    wire NET_304;
    wire NET_305;
    wire NET_306;
    wire NET_307;
    wire NET_308;
    wire NET_309;
    wire NET_310;
    wire NET_311;
    wire NET_312;
    wire NET_313;
    wire NET_314;
    input wire R1C;
    input wire RAG_n;
    input wire RBHG_n;
    input wire RCG_n;
    input wire RGG_n;
    input wire RLG_n;
    input wire RQG_n;
    input wire RUG_n;
    input wire RULOG_n;
    input wire RZG_n;
    input wire SA13;
    input wire SA14;
    input wire SA16;
    output wire SUMA15_n;
    output wire SUMA16_n;
    output wire SUMB15_n;
    output wire SUMB16_n;
    input wire US2SG;
    input wire VCC;
    input wire WAG_n;
    input wire WALSG_n;
    input wire WBG_n;
    input wire WG1G_n;
    input wire WG2G_n;
    input wire WG3G_n;
    input wire WG4G_n;
    input wire WG5G_n;
    input wire WHOMPA;
    input wire WL01_n;
    input wire WL02_n;
    input wire WL12_n;
    output wire WL13_n;
    output wire WL14_n;
    output wire WL15;
    output wire WL15_n;
    output wire WL16;
    output wire WL16_n;
    input wire WLG_n;
    input wire WQG_n;
    input wire WYDG_n;
    input wire WYHIG_n;
    input wire WZG_n;
    input wire XUY01_n;
    input wire XUY02_n;
    output wire XUY13_n;
    output wire XUY14_n;
    wire __A11_1__X1;
    wire __A11_1__X1_n;
    wire __A11_1__X2;
    wire __A11_1__X2_n;
    wire __A11_1__Y1;
    wire __A11_1__Y1_n;
    wire __A11_1__Y2;
    wire __A11_1__Y2_n;
    wire __A11_1___A1_n;
    wire __A11_1___A2_n;
    wire __A11_1___B1_n;
    wire __A11_1___B2_n;
    wire __A11_1___CI_INTERNAL;
    wire __A11_1___G1;
    wire __A11_1___G2;
    wire __A11_1___GEM1;
    wire __A11_1___GEM2;
    wire __A11_1___L1_n;
    wire __A11_1___L2_n;
    wire __A11_1___MWL1;
    wire __A11_1___MWL2;
    wire __A11_1___Q1_n;
    wire __A11_1___Q2_n;
    wire __A11_1___RL1_n;
    wire __A11_1___RL2_n;
    wire __A11_1___RL_OUT_1;
    wire __A11_1___RL_OUT_2;
    wire __A11_1___SUMA1;
    wire __A11_1___SUMA2;
    wire __A11_1___SUMB1;
    wire __A11_1___SUMB2;
    wire __A11_1___WL1;
    wire __A11_1___WL2;
    wire __A11_1___Z1_n;
    wire __A11_1___Z2_n;
    wire __A11_2__X1;
    wire __A11_2__X1_n;
    wire __A11_2__X2;
    wire __A11_2__X2_n;
    wire __A11_2__Y1;
    wire __A11_2__Y1_n;
    wire __A11_2__Y2;
    wire __A11_2__Y2_n;
    wire __A11_2___A1_n;
    wire __A11_2___A2_n;
    wire __A11_2___B1_n;
    wire __A11_2___B2_n;
    wire __A11_2___CI_IN;
    wire __A11_2___CI_INTERNAL;
    wire __A11_2___CO_IN;
    wire __A11_2___CO_OUT;
    wire __A11_2___G1;
    wire __A11_2___G2;
    wire __A11_2___G2_n;
    wire __A11_2___GEM1;
    wire __A11_2___GEM2;
    wire __A11_2___L2_n;
    wire __A11_2___MWL1;
    wire __A11_2___MWL2;
    wire __A11_2___Q1_n;
    wire __A11_2___Q2_n;
    wire __A11_2___RL1_n;
    wire __A11_2___RL2_n;
    wire __A11_2___RL_OUT_1;
    wire __A11_2___RL_OUT_2;
    wire __A11_2___XUY1;
    wire __A11_2___XUY2;
    wire __A11_2___Z1_n;
    wire __A11_2___Z2_n;

    pullup R11001(__A11_2___CO_IN);
    pullup R11002(__A11_1___RL1_n);
    pullup R11003(__A11_1___L1_n);
    pullup R11005(__A11_1___Z1_n);
    pullup R11006(G13_n);
    pullup R11007(__A11_1___RL2_n);
    pullup R11008(__A11_1___L2_n);
    pullup R11009(__A11_1___Z2_n);
    pullup R11010(G14_n);
    pullup R11011(__A11_2___CO_OUT);
    pullup R11012(__A11_2___RL1_n);
    pullup R11013(L15_n);
    pullup R11015(__A11_2___Z1_n);
    pullup R11016(G15_n);
    pullup R11017(__A11_2___RL2_n);
    pullup R11018(__A11_2___L2_n);
    pullup R11019(__A11_2___Z2_n);
    pullup R11020(__A11_2___G2_n);
    U74HC02 U11001(NET_197, A2XG_n, __A11_1___A1_n, NET_192, WYHIG_n, WL13_n, GND, WL12_n, WYDG_n, NET_191, __A11_1__Y1_n, CUG, __A11_1__Y1, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U11002(MONEX, NET_197, __A11_1__X1_n, CLXC, CUG, __A11_1__X1, GND, __A11_1__Y1_n, NET_192, NET_191, __A11_1__Y1, __A11_1__X1_n, __A11_1__X1, VCC, SIM_RST);
    U74HC02 U11003(NET_201, __A11_1__X1_n, __A11_1__Y1_n, XUY13_n, __A11_1__X1, __A11_1__Y1, GND, NET_201, XUY13_n, NET_199, NET_201, __A11_1___SUMA1, __A11_1___CI_INTERNAL, VCC, SIM_RST);
    wire U11004_1_NC;
    wire U11004_2_NC;
    wire U11004_12_NC;
    wire U11004_13_NC;
    U74HC27 U11004(U11004_1_NC, U11004_2_NC, __A11_1___SUMA1, __A11_1___SUMB1, RULOG_n, NET_179, GND, NET_183, __A11_2___XUY1, XUY13_n, CI13_n, U11004_12_NC, U11004_13_NC, VCC, SIM_RST);
    U74HC04 U11005(CI13_n, NET_198, G13_n, __A11_1___GEM1, __A11_1___RL1_n, __A11_1___WL1, GND, WL13_n, __A11_1___WL1, __A11_1___MWL1, __A11_1___RL1_n, NET_149, __A11_1___CI_INTERNAL, VCC, SIM_RST);
    U74HC02 U11006(__A11_1___SUMB1, NET_199, NET_198, NET_182, WAG_n, WL13_n, GND, WL15_n, WALSG_n, NET_184, __A11_1___A1_n, CAG, NET_180, VCC, SIM_RST);
    U74LVC07 U11007(NET_183, __A11_2___CO_IN, NET_177, __A11_1___RL1_n, NET_190, __A11_1___L1_n, GND, __A11_1___Z1_n, NET_213, __A11_1___RL1_n, NET_214, __A11_1___RL1_n, NET_212, VCC, SIM_RST);
    U74HC02 U11008(NET_178, RAG_n, __A11_1___A1_n, NET_181, WLG_n, WL13_n, GND, WL01_n, WALSG_n, NET_188, __A11_1___L1_n, CLG1G, NET_189, VCC, SIM_RST);
    wire U11009_1_NC;
    wire U11009_2_NC;
    wire U11009_3_NC;
    U74HC02 #(0, 0, 1, 0) U11009(U11009_1_NC, U11009_2_NC, U11009_3_NC, NET_186, WQG_n, WL13_n, GND, NET_186, NET_185, __A11_1___Q1_n, __A11_1___Q1_n, CQG, NET_185, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U11010(NET_187, RQG_n, __A11_1___Q1_n, NET_216, WZG_n, WL13_n, GND, NET_216, NET_215, NET_213, __A11_1___Z1_n, CZG, NET_215, VCC, SIM_RST);
    U74HC27 U11011(__A11_1___RL_OUT_1, NET_187, MDT13, R1C, GND, NET_212, GND, NET_219, NET_217, NET_218, NET_204, NET_214, NET_211, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U11012(NET_211, RZG_n, __A11_1___Z1_n, NET_220, WBG_n, WL13_n, GND, NET_220, NET_221, __A11_1___B1_n, __A11_1___B1_n, CBG, NET_221, VCC, SIM_RST);
    U74LVC07 U11013(NET_162, __A11_2___CO_IN, NET_219, __A11_1___RL1_n, NET_203, G13_n, GND, G13_n, NET_202, __A11_1___RL2_n, NET_129, __A11_1___L2_n, NET_139, VCC, SIM_RST);
    U74HC02 U11014(NET_217, RBHG_n, __A11_1___B1_n, NET_218, NET_221, RCG_n, GND, WL12_n, WG3G_n, NET_208, WL14_n, WG4G_n, NET_207, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U11015(NET_182, NET_184, NET_179, NET_178, CH13, NET_177, GND, NET_190, NET_181, NET_188, NET_189, __A11_1___A1_n, NET_180, VCC, SIM_RST);
    U74HC02 U11016(NET_206, L2GDG_n, L12_n, NET_205, WG1G_n, WL13_n, GND, G13_n, CGG, __A11_1___G1, RGG_n, G13_n, NET_204, VCC, SIM_RST);
    U74HC27 #(1, 0, 0) U11017(NET_206, NET_205, GND, __A11_2___XUY2, XUY14_n, NET_162, GND, __A11_1___RL_OUT_1, RLG_n, __A11_1___L1_n, GND, NET_202, __A11_1___G1, VCC, SIM_RST);
    U74HC4002 U11018(NET_203, GND, SA13, NET_208, NET_207, NET_210, GND, NET_209, GND, SA14, NET_156, NET_155, NET_154, VCC, SIM_RST);
    U74HC02 U11019(NET_150, A2XG_n, __A11_1___A2_n, NET_152, WYHIG_n, WL14_n, GND, WL13_n, WYDG_n, NET_151, __A11_1__Y2_n, CUG, __A11_1__Y2, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U11020(MONEX, NET_150, __A11_1__X2_n, CLXC, CUG, __A11_1__X2, GND, __A11_1__Y2_n, NET_152, NET_151, __A11_1__Y2, __A11_1__X2_n, __A11_1__X2, VCC, SIM_RST);
    wire U11021_8_NC;
    wire U11021_9_NC;
    wire U11021_10_NC;
    U74HC02 U11021(NET_144, __A11_1__X2_n, __A11_1__Y2_n, XUY14_n, __A11_1__X2, __A11_1__Y2, GND, U11021_8_NC, U11021_9_NC, U11021_10_NC, NET_144, XUY14_n, NET_147, VCC, SIM_RST);
    wire U11022_1_NC;
    wire U11022_2_NC;
    wire U11022_12_NC;
    wire U11022_13_NC;
    U74HC27 U11022(U11022_1_NC, U11022_2_NC, NET_144, __A11_1___SUMA2, CO14, __A11_2___CI_IN, GND, NET_148, __A11_1___SUMA2, __A11_1___SUMB2, RULOG_n, U11022_12_NC, U11022_13_NC, VCC, SIM_RST);
    U74HC02 U11023(__A11_1___SUMB2, NET_147, NET_149, NET_133, WAG_n, WL14_n, GND, WL16_n, WALSG_n, NET_132, __A11_1___A2_n, CAG, NET_131, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U11024(NET_133, NET_132, NET_148, NET_134, CH14, NET_129, GND, NET_139, NET_167, NET_168, NET_169, __A11_1___A2_n, NET_131, VCC, SIM_RST);
    U74HC02 U11025(NET_134, RAG_n, __A11_1___A2_n, NET_167, WLG_n, WL14_n, GND, WL02_n, WALSG_n, NET_168, __A11_1___L2_n, CLG1G, NET_169, VCC, SIM_RST);
    U74HC27 U11026(RLG_n, __A11_1___L2_n, __A11_1___RL_OUT_2, NET_135, NET_141, NET_140, GND, NET_130, MDT14, R1C, GND, __A11_1___RL_OUT_2, GND, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U11027(NET_171, WQG_n, WL14_n, __A11_1___Q2_n, NET_171, NET_170, GND, __A11_1___Q2_n, CQG, NET_170, RQG_n, __A11_1___Q2_n, NET_135, VCC, SIM_RST);
    U74LVC07 U11028(NET_140, __A11_1___RL2_n, NET_137, __A11_1___Z2_n, NET_130, __A11_1___RL2_n, GND, __A11_1___RL2_n, NET_172, G14_n, NET_154, G14_n, NET_161, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U11029(NET_136, WZG_n, WL14_n, NET_137, NET_136, NET_138, GND, __A11_1___Z2_n, CZG, NET_138, RZG_n, __A11_1___Z2_n, NET_141, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U11030(NET_175, WBG_n, WL14_n, __A11_1___B2_n, NET_175, NET_176, GND, __A11_1___B2_n, CBG, NET_176, RBHG_n, __A11_1___B2_n, NET_174, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U11031(NET_174, NET_173, NET_160, NET_159, __A11_1___G2, NET_161, GND, NET_255, GND, XUY02_n, __A11_2___XUY2, NET_172, NET_153, VCC, SIM_RST);
    U74HC02 U11032(NET_173, NET_176, RCG_n, NET_156, WL13_n, WG3G_n, GND, WL16_n, WG4G_n, NET_155, L2GDG_n, __A11_1___L1_n, NET_160, VCC, SIM_RST);
    wire U11033_11_NC;
    wire U11033_12_NC;
    wire U11033_13_NC;
    U74HC02 U11033(NET_159, WG1G_n, WL14_n, __A11_1___G2, G14_n, CGG, GND, RGG_n, G14_n, NET_153, U11033_11_NC, U11033_12_NC, U11033_13_NC, VCC, SIM_RST);
    wire U11034_10_NC;
    wire U11034_11_NC;
    wire U11034_12_NC;
    wire U11034_13_NC;
    U74HC04 U11034(G14_n, __A11_1___GEM2, __A11_1___RL2_n, __A11_1___WL2, __A11_1___WL2, WL14_n, GND, __A11_1___MWL2, __A11_1___RL2_n, U11034_10_NC, U11034_11_NC, U11034_12_NC, U11034_13_NC, VCC, SIM_RST);
    U74HC02 U11035(NET_290, A2XG_n, __A11_2___A1_n, NET_286, WYHIG_n, WL15_n, GND, WL14_n, WYDG_n, NET_285, __A11_2__Y1_n, CUG, __A11_2__Y1, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U11036(BXVX, NET_290, __A11_2__X1_n, CLXC, CUG, __A11_2__X1, GND, __A11_2__Y1_n, NET_286, NET_285, __A11_2__Y1, __A11_2__X1_n, __A11_2__X1, VCC, SIM_RST);
    U74HC02 U11037(NET_294, __A11_2__X1_n, __A11_2__Y1_n, __A11_2___XUY1, __A11_2__X1, __A11_2__Y1, GND, NET_294, __A11_2___XUY1, NET_291, NET_294, SUMA15_n, __A11_2___CI_INTERNAL, VCC, SIM_RST);
    wire U11038_1_NC;
    wire U11038_2_NC;
    wire U11038_12_NC;
    wire U11038_13_NC;
    U74HC27 U11038(U11038_1_NC, U11038_2_NC, SUMA15_n, SUMB15_n, RULOG_n, NET_272, GND, NET_276, XUY01_n, __A11_2___XUY1, __A11_2___CI_IN, U11038_12_NC, U11038_13_NC, VCC, SIM_RST);
    U74HC04 U11039(__A11_2___CI_IN, NET_292, G15_n, __A11_2___GEM1, __A11_2___RL1_n, WL15, GND, WL15_n, WL15, __A11_2___MWL1, __A11_2___RL1_n, NET_242, __A11_2___CI_INTERNAL, VCC, SIM_RST);
    U74HC02 U11040(SUMB15_n, NET_291, NET_292, NET_275, WAG_n, WL15_n, GND, G16SW_n, WALSG_n, NET_277, __A11_2___A1_n, CAG, NET_273, VCC, SIM_RST);
    U74LVC07 U11041(NET_276, __A11_2___CO_OUT, NET_271, __A11_2___RL1_n, NET_283, L15_n, GND, __A11_2___Z1_n, NET_306, __A11_2___RL1_n, NET_307, __A11_2___RL1_n, NET_305, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U11042(NET_275, NET_277, NET_272, NET_270, CH16, NET_271, GND, NET_283, NET_274, NET_281, NET_282, __A11_2___A1_n, NET_273, VCC, SIM_RST);
    U74HC02 U11043(NET_270, RAG_n, __A11_2___A1_n, NET_274, WLG_n, WL15_n, GND, G01_n, G2LSG_n, NET_281, L15_n, CLG1G, NET_282, VCC, SIM_RST);
    wire U11044_1_NC;
    wire U11044_2_NC;
    wire U11044_3_NC;
    wire U11044_4_NC;
    wire U11044_5_NC;
    wire U11044_6_NC;
    wire U11044_12_NC;
    wire U11044_13_NC;
    U74HC27 U11044(U11044_1_NC, U11044_2_NC, U11044_3_NC, U11044_4_NC, U11044_5_NC, U11044_6_NC, GND, __A11_2___RL_OUT_1, RLG_n, L15_n, VCC, U11044_12_NC, U11044_13_NC, VCC, SIM_RST);
    wire U11045_1_NC;
    wire U11045_2_NC;
    wire U11045_3_NC;
    U74HC02 #(0, 0, 1, 0) U11045(U11045_1_NC, U11045_2_NC, U11045_3_NC, NET_279, WQG_n, WL15_n, GND, NET_279, NET_278, __A11_2___Q1_n, __A11_2___Q1_n, CQG, NET_278, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U11046(NET_280, RQG_n, __A11_2___Q1_n, NET_309, WZG_n, WL15_n, GND, NET_309, NET_308, NET_306, __A11_2___Z1_n, CZG, NET_308, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U11047(NET_304, RZG_n, __A11_2___Z1_n, NET_313, WBG_n, WL15_n, GND, NET_313, NET_314, __A11_2___B1_n, __A11_2___B1_n, CBG, NET_314, VCC, SIM_RST);
    U74HC02 U11048(NET_311, RBHG_n, __A11_2___B1_n, NET_312, NET_314, RCG_n, GND, GND, VCC, NET_301, GND, VCC, NET_300, VCC, SIM_RST);
    U74HC27 U11049(__A11_2___RL_OUT_1, NET_280, MDT15, R1C, __A11_2___RL_OUT_2, NET_305, GND, NET_310, NET_311, NET_312, NET_297, NET_307, NET_304, VCC, SIM_RST);
    U74LVC07 U11050(NET_255, __A11_2___CO_OUT, NET_310, __A11_2___RL1_n, NET_296, G15_n, GND, G15_n, NET_295, __A11_2___RL2_n, NET_222, __A11_2___L2_n, NET_232, VCC, SIM_RST);
    U74HC02 U11051(NET_299, L2GDG_n, __A11_1___L2_n, NET_298, WG1G_n, WL15_n, GND, G15_n, CGG, __A11_2___G1, RGG_n, G15_n, NET_297, VCC, SIM_RST);
    U74HC4002 U11052(NET_296, GND, SA16, NET_301, NET_300, NET_303, GND, NET_302, GND, SA16, NET_249, NET_248, NET_247, VCC, SIM_RST);
    wire U11053_3_NC;
    wire U11053_4_NC;
    wire U11053_5_NC;
    wire U11053_6_NC;
    wire U11053_8_NC;
    wire U11053_9_NC;
    wire U11053_10_NC;
    wire U11053_11_NC;
    U74HC27 #(1, 0, 0) U11053(NET_299, NET_298, U11053_3_NC, U11053_4_NC, U11053_5_NC, U11053_6_NC, GND, U11053_8_NC, U11053_9_NC, U11053_10_NC, U11053_11_NC, NET_295, __A11_2___G1, VCC, SIM_RST);
    U74HC02 U11054(NET_243, A2XG_n, __A11_2___A2_n, NET_245, WYHIG_n, WL16_n, GND, WL16_n, WYDG_n, NET_244, __A11_2__Y2_n, CUG, __A11_2__Y2, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U11055(MONEX, NET_243, __A11_2__X2_n, CLXC, CUG, __A11_2__X2, GND, __A11_2__Y2_n, NET_245, NET_244, __A11_2__Y2, __A11_2__X2_n, __A11_2__X2, VCC, SIM_RST);
    wire U11056_8_NC;
    wire U11056_9_NC;
    wire U11056_10_NC;
    U74HC02 U11056(NET_237, __A11_2__X2_n, __A11_2__Y2_n, __A11_2___XUY2, __A11_2__X2, __A11_2__Y2, GND, U11056_8_NC, U11056_9_NC, U11056_10_NC, NET_237, __A11_2___XUY2, NET_240, VCC, SIM_RST);
    wire U11057_1_NC;
    wire U11057_2_NC;
    wire U11057_12_NC;
    wire U11057_13_NC;
    U74HC27 U11057(U11057_1_NC, U11057_2_NC, NET_237, SUMA16_n, __A11_2___CO_IN, EAC_n, GND, NET_241, SUMA16_n, SUMB16_n, RUG_n, U11057_12_NC, U11057_13_NC, VCC, SIM_RST);
    U74HC02 U11058(SUMB16_n, NET_240, NET_242, NET_226, WAG_n, WL16_n, GND, G16SW_n, WALSG_n, NET_225, __A11_2___A2_n, CAG, NET_224, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U11059(NET_226, NET_225, NET_241, NET_227, CH16, NET_222, GND, NET_232, NET_260, NET_261, NET_262, __A11_2___A2_n, NET_224, VCC, SIM_RST);
    U74HC02 U11060(NET_227, RAG_n, __A11_2___A2_n, NET_260, WLG_n, WL16_n, GND, __A11_2___G2_n, G2LSG_n, NET_261, __A11_2___L2_n, CLG1G, NET_262, VCC, SIM_RST);
    U74HC27 U11061(RLG_n, __A11_2___L2_n, __A11_2___RL_OUT_2, NET_228, NET_234, NET_233, GND, NET_223, MDT16, R1C, US2SG, __A11_2___RL_OUT_2, GND, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U11062(NET_264, WQG_n, WL16_n, __A11_2___Q2_n, NET_264, NET_263, GND, __A11_2___Q2_n, CQG, NET_263, RQG_n, __A11_2___Q2_n, NET_228, VCC, SIM_RST);
    U74LVC07 U11063(NET_233, __A11_2___RL2_n, NET_230, __A11_2___Z2_n, NET_223, __A11_2___RL2_n, GND, __A11_2___RL2_n, NET_265, __A11_2___G2_n, NET_247, __A11_2___G2_n, NET_254, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U11064(NET_229, WZG_n, WL16_n, NET_230, NET_229, NET_231, GND, __A11_2___Z2_n, CZG, NET_231, RZG_n, __A11_2___Z2_n, NET_234, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U11065(NET_268, WBG_n, WL16_n, __A11_2___B2_n, NET_268, NET_269, GND, __A11_2___B2_n, CBG, NET_269, RBHG_n, __A11_2___B2_n, NET_267, VCC, SIM_RST);
    wire U11066_8_NC;
    wire U11066_9_NC;
    wire U11066_10_NC;
    wire U11066_11_NC;
    U74HC27 #(0, 1, 0) U11066(NET_267, NET_266, NET_253, NET_252, __A11_2___G2, NET_254, GND, U11066_8_NC, U11066_9_NC, U11066_10_NC, U11066_11_NC, NET_265, NET_246, VCC, SIM_RST);
    U74HC02 U11067(NET_266, NET_269, RCG_n, NET_249, WL14_n, WG3G_n, GND, WL01_n, WG5G_n, NET_248, L2GDG_n, __A11_2___L2_n, NET_253, VCC, SIM_RST);
    wire U11068_11_NC;
    wire U11068_12_NC;
    wire U11068_13_NC;
    U74HC02 U11068(NET_252, WG2G_n, WL16_n, __A11_2___G2, __A11_2___G2_n, CGG, GND, RGG_n, __A11_2___G2_n, NET_246, U11068_11_NC, U11068_12_NC, U11068_13_NC, VCC, SIM_RST);
    wire U11069_10_NC;
    wire U11069_11_NC;
    wire U11069_12_NC;
    wire U11069_13_NC;
    U74HC04 U11069(__A11_2___G2_n, __A11_2___GEM2, __A11_2___RL2_n, WL16, WL16, WL16_n, GND, __A11_2___MWL2, __A11_2___RL2_n, U11069_10_NC, U11069_11_NC, U11069_12_NC, U11069_13_NC, VCC, SIM_RST);
    U74HC4002 U11070(__A11_1___SUMA1, NET_201, XUY13_n, CI13_n, GND, NET_166, GND, NET_165, NET_144, XUY14_n, __A11_1___CI_INTERNAL, GND, __A11_1___SUMA2, VCC, SIM_RST);
    U74HC4002 U11071(SUMA15_n, NET_294, __A11_2___XUY1, __A11_2___CI_IN, GND, NET_259, GND, NET_258, NET_237, __A11_2___XUY2, __A11_2___CI_INTERNAL, WHOMPA, SUMA16_n, VCC, SIM_RST);
endmodule