`timescale 1ns/1ps
`default_nettype none

module de0_nano_agc(OSC_50, KEY0, EPCS_DATA, EPCS_CSN, EPCS_DCLK, EPCS_ASDI, MT01, MT02, MT03, MT04, MT05, MT06, MT07, MT08, MT09, MT10, MT11, MT12, SNOOP1, SNOOP2);
    input wire OSC_50;
    input wire EPCS_DATA;
    input wire KEY0;
    output wire EPCS_CSN;
    output wire EPCS_DCLK;
    output wire EPCS_ASDI;
    output wire MT01;
    output wire MT02;
    output wire MT03;
    output wire MT04;
    output wire MT05;
    output wire MT06;
    output wire MT07;
    output wire MT08;
    output wire MT09;
    output wire MT10;
    output wire MT11;
    output wire MT12;
     
    output wire SNOOP1;
    output wire SNOOP2;
    
    assign SNOOP1 = EPCS_DCLK;
    assign SNOOP2 = EPCS_ASDI;

    reg VCC = 1;
    reg GND = 0;
    reg SIM_RST = 1;
    reg ALTEST = 0;
    reg BLKUPL_n = 1;
    reg BMGXM = 0;
    reg BMGXP = 0;
    reg BMGYM = 0;
    reg BMGYP = 0;
    reg BMGZM = 0;
    reg BMGZP = 0;
    reg CAURST = 0;
    reg CCH11 = 0;
    reg CCH13 = 0;
    reg CCH14 = 0;
    reg CDUSTB_n = 1;
    reg CDUXD = 0;
    reg CDUXM = 0;
    reg CDUXP = 0;
    reg CDUYD = 0;
    reg CDUYM = 0;
    reg CDUYP = 0;
    reg CDUZD = 0;
    reg CDUZM = 0;
    reg CDUZP = 0;
    reg CH01 = 0;
    reg CH02 = 0;
    reg CH03 = 0;
    reg CH04 = 0;
    reg CH05 = 0;
    reg CH06 = 0;
    reg CH07 = 0;
    reg CH08 = 0;
    reg CH09 = 0;
    reg CH10 = 0;
    reg CH11 = 0;
    reg CH12 = 0;
    reg CH13 = 0;
    reg CH14 = 0;
    reg CH16 = 0;
    reg CHWL01_n = 1;
    reg CHWL02_n = 1;
    reg CHWL03_n = 1;
    reg CHWL04_n = 1;
    reg CHWL05_n = 1;
    reg CHWL06_n = 1;
    reg CHWL07_n = 1;
    reg CHWL08_n = 1;
    reg CHWL09_n = 1;
    reg CHWL10_n = 1;
    reg CHWL11_n = 1;
    reg CHWL12_n = 1;
    reg DBLTEST = 0;
    reg DLKPLS = 0;
    reg E5 = 0;
    reg E6 = 0;
    reg E7_n = 1;
    reg FLTOUT = 0;
    reg GATEX_n = 1;
    reg GATEY_n = 1;
    reg GATEZ_n = 1;
    reg GTONE = 0;
    reg GTSET = 0;
    reg GTSET_n = 1;
    reg HNDRPT = 0;
    reg KYRPT1 = 0;
    reg KYRPT2 = 0;
    reg MAMU = 0;
    reg MDT01 = 0;
    reg MDT02 = 0;
    reg MDT03 = 0;
    reg MDT04 = 0;
    reg MDT05 = 0;
    reg MDT06 = 0;
    reg MDT07 = 0;
    reg MDT08 = 0;
    reg MDT09 = 0;
    reg MDT10 = 0;
    reg MDT11 = 0;
    reg MDT12 = 0;
    reg MDT13 = 0;
    reg MDT14 = 0;
    reg MDT15 = 0;
    reg MDT16 = 0;
    reg MKRPT = 0;
    reg MLDCH = 0;
    reg MLOAD = 0;
    reg MNHNC = 0;
    reg MNHRPT = 0;
    reg MNHSBF = 0;
    reg MONPAR = 0;
    reg MONWBK = 0;
    reg MRDCH = 0;
    reg MREAD = 0;
    reg MSTP = 0;
    reg MSTRT = 0;
    reg MTCSAI = 0;
    reg NHALGA = 0;
    reg NHVFAL = 0;
    reg OVNHRP = 0;
    reg PIPAFL = 0;
    reg PIPPLS_n = 1;
    reg PIPXM = 0;
    reg PIPXP = 0;
    reg PIPYM = 0;
    reg PIPYP = 0;
    reg PIPZM = 0;
    reg PIPZP = 0;
    reg RADRPT = 0;
    reg RCH11_n = 1;
    reg RCH13_n = 1;
    reg RCH14_n = 1;
    reg RCH33_n = 1;
    reg RCHAT_n = 1;
    reg RCHBT_n = 1;
    reg RNRADM = 0;
    reg RNRADP = 0;
    reg SBY = 0;
    reg SCAFAL = 0;
    reg SHAFTD = 0;
    reg SHAFTM = 0;
    reg SHAFTP = 0;
    reg SIGNX = 0;
    reg SIGNY = 0;
    reg SIGNZ = 0;
    reg STNDBY_n = 1;
    reg STRT2 = 0;
    reg T6ON_n = 1;
    reg TEMPIN_n = 1;
    reg TMPOUT = 0;
    reg TRNM = 0;
    reg TRNP = 0;
    reg TRUND = 0;
    reg UPL0 = 0;
    reg UPL1 = 0;
    reg UPRUPT = 0;
    reg VFAIL = 0;
    reg WCH11_n = 1;
    reg WCH13_n = 1;
    reg WCH14_n = 1;
    reg XLNK0 = 0;
    reg XLNK1 = 0;
    reg n2FSFAL = 0;
    wire MGOJAM;

    // Make a 51.2MHz system clock for propagating state, and a 2.048MHz clock
    // that serves as the AGC's clock source
    wire CLOCK;
    wire SYS_CLK;
    pll agc_clock(OSC_50, SYS_CLK, CLOCK);
     
    wire STRT2;
    assign STRT2 = ~KEY0;
     
    fpga_agc AGC(VCC, GND, SIM_RST, SIM_CLK, ALTEST, BLKUPL_n, BMGXM, BMGXP, BMGYM, BMGYP, BMGZM, BMGZP, CAURST, CCH11, CCH13, CCH14, CDUSTB_n, CDUXD, CDUXM, CDUXP, CDUYD, CDUYM, CDUYP, CDUZD, CDUZM, CDUZP, CH01, CH02, CH03, CH04, CH05, CH06, CH07, CH08, CH09, CH10, CH11, CH12, CH13, CH14, CH16, CHWL01_n, CHWL02_n, CHWL03_n, CHWL04_n, CHWL05_n, CHWL06_n, CHWL07_n, CHWL08_n, CHWL09_n, CHWL10_n, CHWL11_n, CHWL12_n, CLOCK, DBLTEST, DLKPLS, E5, E6, E7_n, FLTOUT, GATEX_n, GATEY_n, GATEZ_n, GTONE, GTSET, GTSET_n, HNDRPT, KYRPT1, KYRPT2, MAMU, MDT01, MDT02, MDT03, MDT04, MDT05, MDT06, MDT07, MDT08, MDT09, MDT10, MDT11, MDT12, MDT13, MDT14, MDT15, MDT16, MKRPT, MLDCH, MLOAD, MNHNC, MNHRPT, MNHSBF, MONPAR, MONWBK, MRDCH, MREAD, MSTP, MSTRT, MTCSAI, NHALGA, NHVFAL, OVNHRP, PIPAFL, PIPPLS_n, PIPXM, PIPXP, PIPYM, PIPYP, PIPZM, PIPZP, RADRPT, RCH11_n, RCH13_n, RCH14_n, RCH33_n, RCHAT_n, RCHBT_n, RNRADM, RNRADP, SBY, SCAFAL, SHAFTD, SHAFTM, SHAFTP, SIGNX, SIGNY, SIGNZ, STNDBY_n, STRT2, T6ON_n, TEMPIN_n, TMPOUT, TRNM, TRNP, TRUND, UPL0, UPL1, UPRUPT, VFAIL, WCH11_n, WCH13_n, WCH14_n, XLNK0, XLNK1, n2FSFAL, MGOJAM, MT01, MT02, MT03, MT04, MT05, MT06, MT07, MT08, MT09, MT10, MT11, MT12);

endmodule
