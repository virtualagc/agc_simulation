`timescale 1ns/1ps
`default_nettype none

module memory_timing_addressing(VCC, GND, SIM_RST, SIM_CLK, GOJAM, STRT2, PHS2_n, PHS3_n, PHS4_n, T01, T01_n, T02_n, T03, T03_n, T04_n, T05, T05_n, T06, T06_n, T07, T07_n, T08, T08_n, T09, T10, T10_n, T11, T12_n, T12A, S01, S01_n, S02, S02_n, S03, S03_n, S04, S04_n, S05, S05_n, S06, S06_n, S07, S07_n, S08, S08_n, S09, S09_n, S10_n, S11, S12, EB9, EB10, EB11_n, CHINC, DV3764, GOJ1, INOUT, MP1, TCSAJ3, SCAD, TIMR, MAMU, MNHSBF, STBE, STBF, SBF, STRGAT, TPARG_n, XB0, XB0_n, XB1, XB1_n, XB2, XB2_n, XB3, XB3_n, XB4, XB4_n, XB5, XB5_n, XB6, XB6_n, XB7, XB7_n, XT0_n, XT1_n, XT2_n, XT3_n, XT4_n, XT5_n, XT6_n, YB0_n, YT0_n, SETAB, SETCD, RESETA, RESETB, RESETC, RESETD, CLROPE, IL01, IL02, IL03, IL04, IL05, IL06, IL07, SBE, SETEK, WEX, WEY, ZID, XB7E, XB1E, XB2E, XB3E, XB4E, XB5E, XB6E, XT7E, XT1E, XT2E, XT3E, XT4E, XT5E, XT6E, YB3E, YB1E, YB2E, YT7E, YT1E, YT2E, YT3E, YT4E, YT5E, YT6E);
    input wire VCC;
    input wire GND;
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire CHINC;
    output wire CLROPE;
    input wire DV3764;
    input wire EB10;
    input wire EB11_n;
    input wire EB9;
    input wire GOJ1;
    input wire GOJAM;
    output wire IL01;
    output wire IL02;
    output wire IL03;
    output wire IL04;
    output wire IL05;
    output wire IL06;
    output wire IL07;
    input wire INOUT;
    input wire MAMU;
    input wire MNHSBF;
    input wire MP1;
    input wire PHS2_n;
    input wire PHS3_n;
    input wire PHS4_n;
    output wire RESETA;
    output wire RESETB;
    output wire RESETC;
    output wire RESETD;
    input wire S01;
    input wire S01_n;
    input wire S02;
    input wire S02_n;
    input wire S03;
    input wire S03_n;
    input wire S04;
    input wire S04_n;
    input wire S05;
    input wire S05_n;
    input wire S06;
    input wire S06_n;
    input wire S07;
    input wire S07_n;
    input wire S08;
    input wire S08_n;
    input wire S09;
    input wire S09_n;
    input wire S10_n;
    input wire S11;
    input wire S12;
    output wire SBE;
    output wire SBF;
    input wire SCAD;
    output wire SETAB;
    output wire SETCD;
    output wire SETEK;
    output wire STBE;
    output wire STBF;
    output wire STRGAT;
    input wire STRT2;
    input wire T01;
    input wire T01_n;
    input wire T02_n;
    input wire T03;
    input wire T03_n;
    input wire T04_n;
    input wire T05;
    input wire T05_n;
    input wire T06;
    input wire T06_n;
    input wire T07;
    input wire T07_n;
    input wire T08;
    input wire T08_n;
    input wire T09;
    input wire T10;
    input wire T10_n;
    input wire T11;
    input wire T12A;
    input wire T12_n;
    input wire TCSAJ3;
    input wire TIMR;
    output wire TPARG_n;
    output wire WEX;
    output wire WEY;
    output wire XB0;
    output wire XB0_n;
    output wire XB1;
    output wire XB1E;
    output wire XB1_n;
    output wire XB2;
    output wire XB2E;
    output wire XB2_n;
    output wire XB3;
    output wire XB3E;
    output wire XB3_n;
    output wire XB4;
    output wire XB4E;
    output wire XB4_n;
    output wire XB5;
    output wire XB5E;
    output wire XB5_n;
    output wire XB6;
    output wire XB6E;
    output wire XB6_n;
    output wire XB7;
    output wire XB7E;
    output wire XB7_n;
    output wire XT0_n;
    output wire XT1E;
    output wire XT1_n;
    output wire XT2E;
    output wire XT2_n;
    output wire XT3E;
    output wire XT3_n;
    output wire XT4E;
    output wire XT4_n;
    output wire XT5E;
    output wire XT5_n;
    output wire XT6E;
    output wire XT6_n;
    output wire XT7E;
    output wire YB0_n;
    output wire YB1E;
    output wire YB2E;
    output wire YB3E;
    output wire YT0_n;
    output wire YT1E;
    output wire YT2E;
    output wire YT3E;
    output wire YT4E;
    output wire YT5E;
    output wire YT6E;
    output wire YT7E;
    output wire ZID;
    wire __A14_1__CLEARA;
    wire __A14_1__CLEARB;
    wire __A14_1__CLEARC;
    wire __A14_1__CLEARD;
    wire __A14_1__ERAS; //FPGA#wand
    wire __A14_1__ERAS_n;
    wire __A14_1__FNERAS_n;
    wire __A14_1__IHENV;
    wire __A14_1__REDRST;
    wire __A14_1__REX;
    wire __A14_1__REY;
    wire __A14_1__ROP_n;
    wire __A14_1__RSTKX_n;
    wire __A14_1__RSTKY_n;
    wire __A14_1__RSTK_n;
    wire __A14_1__S08A;
    wire __A14_1__S08A_n;
    wire __A14_1__SBESET;
    wire __A14_1__SBFSET; //FPGA#wand
    wire __A14_1__SETAB_n;
    wire __A14_1__SETCD_n;
    wire __A14_1__TPGE; //FPGA#wand
    wire __A14_1__TPGF; //FPGA#wand
    wire __A14_2__EAD09;
    wire __A14_2__EAD09_n;
    wire __A14_2__EAD10;
    wire __A14_2__EAD10_n;
    wire __A14_2__EAD11;
    wire __A14_2__EAD11_n;
    wire __A14_2__IL01_n;
    wire __A14_2__IL02_n;
    wire __A14_2__IL03_n;
    wire __A14_2__IL04_n;
    wire __A14_2__IL05_n;
    wire __A14_2__IL06_n;
    wire __A14_2__IL07_n;
    wire __A14_2__ILP;
    wire __A14_2__ILP_n;
    wire __A14_2__RILP1;
    wire __A14_2__RILP1_n;
    wire __A14_2__XB0E;
    wire __A14_2__XT0;
    wire __A14_2__XT0E;
    wire __A14_2__XT1;
    wire __A14_2__XT2;
    wire __A14_2__XT3;
    wire __A14_2__XT4;
    wire __A14_2__XT5;
    wire __A14_2__XT6;
    wire __A14_2__XT7;
    wire __A14_2__XT7_n;
    wire __A14_2__YB0;
    wire __A14_2__YB0E;
    wire __A14_2__YB1;
    wire __A14_2__YB1_n;
    wire __A14_2__YB2;
    wire __A14_2__YB2_n;
    wire __A14_2__YB3;
    wire __A14_2__YB3_n;
    wire __A14_2__YT0;
    wire __A14_2__YT0E;
    wire __A14_2__YT1;
    wire __A14_2__YT1_n;
    wire __A14_2__YT2;
    wire __A14_2__YT2_n;
    wire __A14_2__YT3;
    wire __A14_2__YT3_n;
    wire __A14_2__YT4;
    wire __A14_2__YT4_n;
    wire __A14_2__YT5;
    wire __A14_2__YT5_n;
    wire __A14_2__YT6;
    wire __A14_2__YT6_n;
    wire __A14_2__YT7;
    wire __A14_2__YT7_n;
    wire __A14_NET_192;
    wire __A14_NET_194;
    wire __A14_NET_196;
    wire __A14_NET_198;
    wire __A14_NET_199;
    wire __A14_NET_200;
    wire __A14_NET_202;
    wire __A14_NET_203;
    wire __A14_NET_204;
    wire __A14_NET_205;
    wire __A14_NET_206;
    wire __A14_NET_207;
    wire __A14_NET_208;
    wire __A14_NET_209;
    wire __A14_NET_210;
    wire __A14_NET_211;
    wire __A14_NET_212;
    wire __A14_NET_213;
    wire __A14_NET_214;
    wire __A14_NET_215;
    wire __A14_NET_216;
    wire __A14_NET_217;
    wire __A14_NET_218;
    wire __A14_NET_219;
    wire __A14_NET_220;
    wire __A14_NET_221;
    wire __A14_NET_222;
    wire __A14_NET_223;
    wire __A14_NET_224;
    wire __A14_NET_225;
    wire __A14_NET_226;
    wire __A14_NET_231;
    wire __A14_NET_232;
    wire __A14_NET_233;
    wire __A14_NET_234;
    wire __A14_NET_235;
    wire __A14_NET_236;
    wire __A14_NET_237;
    wire __A14_NET_238;
    wire __A14_NET_239;
    wire __A14_NET_240;
    wire __A14_NET_241;
    wire __A14_NET_242;
    wire __A14_NET_246;
    wire __A14_NET_247;
    wire __A14_NET_248;
    wire __A14_NET_249;
    wire __A14_NET_250;
    wire __A14_NET_251;
    wire __A14_NET_252;
    wire __A14_NET_253;
    wire __A14_NET_254;
    wire __A14_NET_255;
    wire __A14_NET_256;
    wire __A14_NET_257;
    wire __A14_NET_258;
    wire __A14_NET_259;
    wire __A14_NET_260;
    wire __A14_NET_261;
    wire __A14_NET_262;
    wire __A14_NET_263;
    wire __A14_NET_264;
    wire __A14_NET_265;
    wire __A14_NET_266;
    wire __A14_NET_267;
    wire __A14_NET_268;
    wire __A14_NET_269;
    wire __A14_NET_270;
    wire __A14_NET_271;
    wire __A14_NET_272;
    wire __A14_NET_274;
    wire __A14_NET_275;
    wire __A14_NET_276;
    wire __A14_NET_279;
    wire __A14_NET_280;
    wire __A14_NET_285;
    wire __A14_NET_286;
    wire __A14_NET_287;
    wire __A14_NET_288;
    wire __A14_NET_289;
    wire __A14_NET_290;
    wire __A14_NET_292;
    wire __A14_NET_295;
    wire __A14_NET_296;
    wire __A14_NET_297;
    wire __A14_NET_300;
    wire __A14_NET_301;
    wire __A14_NET_306;
    wire __A14_NET_308;

    pullup R14001(__A14_1__SBFSET);
    pullup R14002(__A14_1__TPGF);
    pullup R14003(__A14_1__ERAS);
    pullup R14004(__A14_1__TPGE);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b1) U14001(__A14_1__ROP_n, S11, S12, __A14_NET_210, T08_n, PHS3_n, GND, __A14_NET_210, __A14_NET_211, __A14_NET_209, __A14_NET_212, __A14_NET_213, __A14_NET_206, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14002(__A14_NET_209, T09, __A14_1__ROP_n, __A14_NET_209, T08, __A14_NET_212, GND, __A14_NET_213, __A14_NET_206, __A14_NET_207, TIMR, __A14_NET_211, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14003(T01_n, __A14_NET_207, __A14_NET_206, __A14_1__IHENV, __A14_NET_219, __A14_1__SETAB_n, GND, SETAB, __A14_1__SETAB_n, __A14_1__SETCD_n, __A14_NET_220, SETCD, __A14_1__SETCD_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14004(TIMR, __A14_NET_207, PHS4_n, __A14_1__ROP_n, T10_n, __A14_NET_208, GND, __A14_NET_214, T05_n, PHS3_n, __A14_1__ROP_n, __A14_NET_205, __A14_NET_218, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U14005(__A14_NET_218, __A14_NET_205, __A14_NET_208, __A14_NET_219, S09, __A14_NET_218, GND, __A14_NET_218, S09_n, __A14_NET_220, __A14_NET_214, __A14_NET_215, __A14_NET_199, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14006(__A14_NET_199, T08, __A14_NET_199, S09, S08, __A14_NET_216, GND, __A14_NET_196, __A14_NET_199, S09, S08_n, __A14_NET_215, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74HC02 U14007(__A14_NET_217, __A14_1__CLEARA, __A14_NET_216, __A14_NET_198, __A14_1__CLEARB, __A14_NET_196, GND, __A14_1__CLEARC, __A14_NET_200, __A14_NET_202, __A14_1__CLEARD, __A14_NET_194, __A14_NET_192, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14008(__A14_NET_217, RESETA, __A14_NET_198, RESETB, __A14_NET_202, RESETC, GND, RESETD, __A14_NET_192, __A14_1__S08A_n, S08, __A14_1__S08A, S08_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14009(__A14_NET_199, S08, __A14_NET_199, S09_n, S08_n, __A14_NET_194, GND, STBF, GOJAM, __A14_NET_204, __A14_NET_203, __A14_NET_200, S09_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U14010(__A14_1__CLEARA, __A14_1__SETAB_n, __A14_1__S08A_n, __A14_1__CLEARB, __A14_1__SETAB_n, __A14_1__S08A, GND, __A14_1__SETCD_n, __A14_1__S08A_n, __A14_1__CLEARC, __A14_1__SETCD_n, __A14_1__S08A, __A14_1__CLEARD, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U14011(__A14_NET_203, STBF, __A14_1__SBFSET, __A14_NET_204, T07_n, PHS3_n, GND, T02_n, __A14_1__ROP_n, __A14_NET_235, __A14_NET_235, STRGAT, __A14_NET_236, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14012(__A14_NET_203, SBF, __A14_1__ROP_n, __A14_NET_260, S07_n, __A14_2__IL07_n, GND, WEX, __A14_NET_250, WEY, __A14_NET_249, __A14_1__ERAS_n, __A14_1__ERAS, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14013(MNHSBF, MP1, __A14_1__ROP_n, T05_n, DV3764, __A14_NET_280, GND, STRGAT, __A14_NET_236, T08, GOJAM, __A14_NET_279, PHS4_n, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U14014(__A14_NET_279, __A14_1__SBFSET, __A14_NET_280, __A14_1__SBFSET, __A14_NET_285, __A14_1__TPGF, GND, __A14_1__TPGF, __A14_NET_286, __A14_1__ERAS, __A14_NET_231, __A14_1__ERAS, __A14_NET_226, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC4002 U14015(__A14_NET_285, __A14_1__ROP_n, T08_n, DV3764, GOJ1,  , GND,  , GOJAM, TCSAJ3, PHS2_n, MP1, __A14_NET_286, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14016(T02_n, __A14_NET_260, __A14_NET_265, T03, GOJAM, __A14_NET_258, GND, __A14_NET_263, __A14_NET_262, T07, GOJAM, __A14_NET_264, __A14_NET_265, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U14017(__A14_NET_259, __A14_1__ROP_n, T10_n, __A14_NET_265, __A14_NET_259, __A14_NET_258, GND, __A14_NET_264, __A14_NET_263, __A14_NET_262, T01, __A14_NET_261, __A14_NET_253, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U14018(__A14_NET_261, __A14_NET_253, __A14_NET_252, __A14_NET_252, T12_n, PHS3_n, GND, T12A, __A14_NET_261, __A14_NET_257, __A14_NET_251, __A14_NET_255, __A14_NET_250, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14019(__A14_NET_257, TIMR, __A14_NET_257, TIMR, __A14_NET_249, __A14_NET_248, GND, __A14_NET_254, TIMR, T11, __A14_NET_256, __A14_NET_251, __A14_NET_250, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b0, 1'b0) U14020(__A14_NET_249, __A14_NET_248, __A14_NET_276, __A14_NET_256, __A14_NET_254, __A14_NET_270, GND, __A14_NET_256, T10, __A14_NET_255, T05_n, __A14_1__ERAS_n, __A14_NET_275, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14021(__A14_NET_242, __A14_NET_224, __A14_1__ERAS_n, PHS3_n, T03_n, __A14_NET_223, GND, __A14_NET_274, __A14_1__FNERAS_n, T12A, GOJAM, __A14_NET_232, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U14022(__A14_1__FNERAS_n, __A14_NET_275, __A14_NET_274, __A14_NET_271, __A14_1__FNERAS_n, T10_n, GND, __A14_NET_266, __A14_NET_270, __A14_NET_269, T02_n, PHS4_n, __A14_NET_268, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14023(T10_n, __A14_1__FNERAS_n, __A14_1__FNERAS_n, T10_n, PHS3_n, __A14_NET_270, GND, __A14_NET_266, TIMR, __A14_NET_268, __A14_NET_269, __A14_NET_276, PHS4_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14024(TIMR, T01, __A14_NET_222, GOJAM, __A14_1__REDRST, __A14_NET_221, GND, __A14_NET_225, __A14_NET_233, GOJAM, __A14_1__REDRST, __A14_NET_272, __A14_NET_267, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U14025(__A14_NET_267, __A14_NET_272, __A14_NET_271, ZID, __A14_NET_267, STRT2, GND, __A14_1__ERAS_n, T03_n, __A14_NET_234, __A14_NET_234, __A14_NET_232, __A14_NET_242, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U14026(__A14_NET_231, TCSAJ3, S11, S12, INOUT,  , GND,  , CHINC, GOJ1, MP1, MAMU, __A14_NET_226, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b1) U14027(SETEK, STRT2, __A14_NET_242, __A14_NET_224, T06_n, PHS3_n, GND, __A14_NET_223, __A14_NET_221, __A14_NET_222, __A14_NET_237, __A14_NET_225, __A14_NET_233, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14028(__A14_NET_222, __A14_1__REY, __A14_NET_233, __A14_1__REX, __A14_NET_239, SBE, GND, __A14_1__RSTK_n, __A14_NET_269, __A14_1__RSTKY_n, __A14_1__RSTK_n, __A14_1__RSTKX_n, __A14_1__RSTK_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14029(__A14_1__ERAS_n, T03_n, GOJAM, T05, __A14_NET_239, STBE, GND, __A14_1__SBESET, T04_n, __A14_1__ERAS_n, SCAD, __A14_NET_237, PHS4_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U14030(__A14_1__REDRST, __A14_NET_238, T05, __A14_NET_238, __A14_NET_241, __A14_NET_240, GND, __A14_NET_238, T06, __A14_NET_240, T05_n, PHS3_n, __A14_NET_241, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U14031(__A14_NET_239, STBE, __A14_1__SBESET, __A14_NET_247, T05_n, PHS3_n, GND, __A14_1__TPGF, __A14_1__TPGE, TPARG_n, S07, S08, __A14_2__YB0, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14032(SCAD, __A14_1__ERAS_n, S01, S02, S03, XB0, GND, XB1, S01_n, S02, S03, __A14_NET_246, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U14033(__A14_NET_246, __A14_1__TPGE, __A14_NET_247, __A14_1__TPGE,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4
    U74HC04 U14034(XB0, XB0_n, XB0_n, __A14_2__XB0E, XB1, XB1_n, GND, XB1E, XB1_n, XB2_n, XB2, XB2E, XB2_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14035(S01, S02_n, S01_n, S02_n, S03, XB3, GND, XB4, S01, S02, S03_n, XB2, S03, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14036(XB3, XB3_n, XB3_n, XB3E, XB4, XB4_n, GND, XB4E, XB4_n, XB5_n, XB5, XB5E, XB5_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14037(S01_n, S02, S01, S02_n, S03_n, XB6, GND, XB7, S01_n, S02_n, S03_n, XB5, S03_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14038(XB6, XB6_n, XB6_n, XB6E, XB7, XB7_n, GND, XB7E, XB7_n, YB0_n, __A14_2__YB0, __A14_2__YB0E, YB0_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U14039(__A14_2__YB1, S07_n, S08, __A14_2__YB2, S07, S08_n, GND, S07_n, S08_n, __A14_2__YB3, EB9, S10_n, __A14_NET_287, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14040(__A14_2__YB1, __A14_2__YB1_n, __A14_2__YB1_n, YB1E, __A14_2__YB2, __A14_2__YB2_n, GND, YB2E, __A14_2__YB2_n, __A14_2__YB3_n, __A14_2__YB3, YB3E, __A14_2__YB3_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14041(S04, S05, S04_n, S05, S06, __A14_2__XT1, GND, __A14_2__XT2, S04, S05_n, S06, __A14_2__XT0, S06, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14042(__A14_2__XT0, XT0_n, XT0_n, __A14_2__XT0E, __A14_2__XT1, XT1_n, GND, XT1E, XT1_n, XT2_n, __A14_2__XT2, XT2E, XT2_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14043(S04_n, S05_n, S04, S05, S06_n, __A14_2__XT4, GND, __A14_2__XT5, S04_n, S05, S06_n, __A14_2__XT3, S06, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14044(__A14_2__XT3, XT3_n, XT3_n, XT3E, __A14_2__XT4, XT4_n, GND, XT4E, XT4_n, XT5_n, __A14_2__XT5, XT5E, XT5_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14045(S04, S05_n, S04_n, S05_n, S06_n, __A14_2__XT7, GND, __A14_2__EAD11, S09_n, S10_n, EB11_n, __A14_2__XT6, S06_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14046(__A14_2__XT6, XT6_n, XT6_n, XT6E, __A14_2__XT7, __A14_2__XT7_n, GND, XT7E, __A14_2__XT7_n, __A14_2__EAD09_n, __A14_2__EAD09, __A14_2__EAD10_n, __A14_2__EAD10, VCC, SIM_RST, SIM_CLK);
    U74HC02 U14047(__A14_2__EAD09, __A14_NET_287, S09_n, __A14_NET_306, EB10, S09_n, GND, S10_n, __A14_NET_306, __A14_2__EAD10, __A14_2__YB0, __A14_2__YB3, __A14_2__RILP1, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14048(__A14_2__EAD11, __A14_2__EAD11_n, __A14_2__YT0, YT0_n, YT0_n, __A14_2__YT0E, GND, __A14_2__YT1_n, __A14_2__YT1, YT1E, __A14_2__YT1_n, __A14_2__YT2_n, __A14_2__YT2, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14049(__A14_2__EAD09, __A14_2__EAD10, __A14_2__EAD09_n, __A14_2__EAD10, __A14_2__EAD11, __A14_2__YT1, GND, __A14_2__YT2, __A14_2__EAD09, __A14_2__EAD10_n, __A14_2__EAD11, __A14_2__YT0, __A14_2__EAD11, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14050(__A14_2__YT2_n, YT2E, __A14_2__YT3, __A14_2__YT3_n, __A14_2__YT3_n, YT3E, GND, __A14_2__YT4_n, __A14_2__YT4, YT4E, __A14_2__YT4_n, __A14_2__YT5_n, __A14_2__YT5, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14051(__A14_2__EAD09_n, __A14_2__EAD10_n, __A14_2__EAD09, __A14_2__EAD10, __A14_2__EAD11_n, __A14_2__YT4, GND, __A14_2__YT5, __A14_2__EAD09_n, __A14_2__EAD10, __A14_2__EAD11_n, __A14_2__YT3, __A14_2__EAD11, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14052(__A14_2__YT5_n, YT5E, __A14_2__YT6, __A14_2__YT6_n, __A14_2__YT6_n, YT6E, GND, __A14_2__YT7_n, __A14_2__YT7, YT7E, __A14_2__YT7_n, __A14_NET_288, __A14_NET_292, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14053(__A14_2__EAD09, __A14_2__EAD10_n, __A14_2__EAD09_n, __A14_2__EAD10_n, __A14_2__EAD11_n, __A14_2__YT7, GND, __A14_NET_290, __A14_NET_292, __A14_2__RILP1, __A14_NET_289, __A14_2__YT6, __A14_2__EAD11_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U14054(__A14_NET_292, XB0, XB3, XB5, XB6,  , GND,  , __A14_2__XT0, __A14_2__XT3, __A14_2__XT5, __A14_2__XT6, __A14_NET_289, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14055(__A14_NET_289, __A14_NET_308, __A14_2__RILP1, __A14_2__RILP1_n, __A14_NET_300, __A14_NET_301, GND, __A14_2__ILP_n, __A14_NET_300, __A14_2__ILP, __A14_NET_301, IL01, S01, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14056(__A14_NET_288, __A14_2__RILP1, __A14_NET_288, __A14_2__RILP1_n, __A14_NET_289, __A14_NET_297, GND, __A14_NET_296, __A14_NET_292, __A14_2__RILP1_n, __A14_NET_308, __A14_NET_295, __A14_NET_308, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U14057(__A14_NET_300, __A14_NET_290, __A14_NET_295, __A14_NET_297, __A14_NET_296,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U14058(S01_n, __A14_2__IL01_n, S02, IL02, S02_n, __A14_2__IL02_n, GND, IL03, S03, __A14_2__IL03_n, S03_n, IL04, S04, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14059(S04_n, __A14_2__IL04_n, S05, IL05, S05_n, __A14_2__IL05_n, GND, IL06, S06, __A14_2__IL06_n, S06_n, IL07, S07, VCC, SIM_RST, SIM_CLK);
    U74HC02 U14060(CLROPE, STRT2, __A14_NET_262,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
endmodule