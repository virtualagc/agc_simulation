`timescale 1ns/1ps
`default_nettype none

module four_bit_1(VCC, GND, SIM_RST, SIM_CLK, A2XG_n, CAG, CBG, CGG, CLG1G, CLXC, CQG, CUG, CZG, L2GDG_n, RAG_n, RCG_n, RGG_n, RLG_n, RQG_n, RZG_n, WAG_n, WALSG_n, WBG_n, WLG_n, WQG_n, WZG_n, CI01_n, MONEX, PONEX, TWOX, XUY05_n, XUY06_n, CH01, CH02, CH03, CH04, G01ED, G02ED, G03ED, G04ED, MCRO_n, G2LSG_n, G05_n, G06_n, G07_n, MDT01, MDT02, MDT03, MDT04, SA01, SA02, SA03, SA04, RBLG_n, RULOG_n, WL05_n, WL06_n, WG1G_n, WG3G_n, WG4G_n, WYDLOG_n, WYDG_n, WYLOG_n, RB1, R1C, R15, RB2, WL16_n, WHOMP, WHOMPA, CI05_n, CO06, G01, G01_n, G02, G03, G04, L01_n, L02_n, L04_n, RL01_n, RL02_n, RL03_n, RL04_n, SUMA01_n, SUMB01_n, SUMA02_n, SUMB02_n, SUMA03_n, SUMB03_n, WL01, WL01_n, WL02, WL02_n, WL03, WL03_n, WL04, WL04_n, XUY01_n, XUY02_n, GEM01, GEM02, GEM03, GEM04);
    input wire VCC;
    input wire GND;
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire A2XG_n;
    input wire CAG;
    input wire CBG;
    input wire CGG;
    input wire CH01;
    input wire CH02;
    input wire CH03;
    input wire CH04;
    input wire CI01_n;
    output wire CI05_n;
    input wire CLG1G;
    input wire CLXC;
    output wire CO06; //FPGA#wand
    input wire CQG;
    input wire CUG;
    input wire CZG;
    output wire G01;
    input wire G01ED;
    inout wire G01_n; //FPGA#wand
    output wire G02;
    input wire G02ED;
    output wire G03;
    input wire G03ED;
    output wire G04;
    input wire G04ED;
    input wire G05_n;
    input wire G06_n;
    input wire G07_n;
    input wire G2LSG_n;
    output wire GEM01;
    output wire GEM02;
    output wire GEM03;
    output wire GEM04;
    inout wire L01_n; //FPGA#wand
    inout wire L02_n; //FPGA#wand
    inout wire L04_n; //FPGA#wand
    input wire L2GDG_n;
    input wire MCRO_n;
    input wire MDT01;
    input wire MDT02;
    input wire MDT03;
    input wire MDT04;
    input wire MONEX;
    input wire PONEX;
    input wire R15;
    input wire R1C;
    input wire RAG_n;
    input wire RB1;
    input wire RB2;
    input wire RBLG_n;
    input wire RCG_n;
    input wire RGG_n;
    inout wire RL01_n; //FPGA#wand
    inout wire RL02_n; //FPGA#wand
    inout wire RL03_n; //FPGA#wand
    inout wire RL04_n; //FPGA#wand
    input wire RLG_n;
    input wire RQG_n;
    input wire RULOG_n;
    input wire RZG_n;
    input wire SA01;
    input wire SA02;
    input wire SA03;
    input wire SA04;
    output wire SUMA01_n;
    output wire SUMA02_n;
    output wire SUMA03_n;
    output wire SUMB01_n;
    output wire SUMB02_n;
    output wire SUMB03_n;
    input wire TWOX;
    input wire WAG_n;
    input wire WALSG_n;
    input wire WBG_n;
    input wire WG1G_n;
    input wire WG3G_n;
    input wire WG4G_n;
    input wire WHOMP;
    input wire WHOMPA;
    output wire WL01;
    output wire WL01_n;
    output wire WL02;
    output wire WL02_n;
    output wire WL03;
    output wire WL03_n;
    output wire WL04;
    output wire WL04_n;
    input wire WL05_n;
    input wire WL06_n;
    input wire WL16_n;
    input wire WLG_n;
    input wire WQG_n;
    input wire WYDG_n;
    input wire WYDLOG_n;
    input wire WYLOG_n;
    input wire WZG_n;
    output wire XUY01_n;
    output wire XUY02_n;
    input wire XUY05_n;
    input wire XUY06_n;
    wire __A08_1__X1;
    wire __A08_1__X1_n;
    wire __A08_1__X2;
    wire __A08_1__X2_n;
    wire __A08_1__Y1;
    wire __A08_1__Y1_n;
    wire __A08_1__Y2;
    wire __A08_1__Y2_n;
    wire __A08_1___A1_n;
    wire __A08_1___A2_n;
    wire __A08_1___B1_n;
    wire __A08_1___B2_n;
    wire __A08_1___CI_INTERNAL;
    wire __A08_1___G2_n; //FPGA#wand
    wire __A08_1___MWL1;
    wire __A08_1___MWL2;
    wire __A08_1___Q1_n;
    wire __A08_1___Q2_n;
    wire __A08_1___RL_OUT_1;
    wire __A08_1___RL_OUT_2;
    wire __A08_1___Z1_n; //FPGA#wand
    wire __A08_1___Z2_n; //FPGA#wand
    wire __A08_2__X1;
    wire __A08_2__X1_n;
    wire __A08_2__X2;
    wire __A08_2__X2_n;
    wire __A08_2__Y1;
    wire __A08_2__Y1_n;
    wire __A08_2__Y2;
    wire __A08_2__Y2_n;
    wire __A08_2___A1_n;
    wire __A08_2___A2_n;
    wire __A08_2___B1_n;
    wire __A08_2___B2_n;
    wire __A08_2___CI_IN;
    wire __A08_2___CI_INTERNAL;
    wire __A08_2___CO_IN; //FPGA#wand
    wire __A08_2___G1_n; //FPGA#wand
    wire __A08_2___G2_n; //FPGA#wand
    wire __A08_2___L1_n; //FPGA#wand
    wire __A08_2___MWL1;
    wire __A08_2___MWL2;
    wire __A08_2___Q1_n;
    wire __A08_2___Q2_n;
    wire __A08_2___RL_OUT_1;
    wire __A08_2___RL_OUT_2;
    wire __A08_2___SUMA2;
    wire __A08_2___SUMB2;
    wire __A08_2___XUY1;
    wire __A08_2___XUY2;
    wire __A08_2___Z1_n; //FPGA#wand
    wire __A08_2___Z2_n; //FPGA#wand
    wire __A08_NET_137;
    wire __A08_NET_138;
    wire __A08_NET_139;
    wire __A08_NET_140;
    wire __A08_NET_141;
    wire __A08_NET_142;
    wire __A08_NET_143;
    wire __A08_NET_144;
    wire __A08_NET_145;
    wire __A08_NET_146;
    wire __A08_NET_147;
    wire __A08_NET_148;
    wire __A08_NET_149;
    wire __A08_NET_152;
    wire __A08_NET_155;
    wire __A08_NET_156;
    wire __A08_NET_157;
    wire __A08_NET_158;
    wire __A08_NET_159;
    wire __A08_NET_160;
    wire __A08_NET_161;
    wire __A08_NET_162;
    wire __A08_NET_163;
    wire __A08_NET_164;
    wire __A08_NET_167;
    wire __A08_NET_168;
    wire __A08_NET_169;
    wire __A08_NET_170;
    wire __A08_NET_175;
    wire __A08_NET_176;
    wire __A08_NET_177;
    wire __A08_NET_178;
    wire __A08_NET_179;
    wire __A08_NET_180;
    wire __A08_NET_181;
    wire __A08_NET_182;
    wire __A08_NET_183;
    wire __A08_NET_184;
    wire __A08_NET_185;
    wire __A08_NET_186;
    wire __A08_NET_187;
    wire __A08_NET_188;
    wire __A08_NET_189;
    wire __A08_NET_190;
    wire __A08_NET_191;
    wire __A08_NET_192;
    wire __A08_NET_193;
    wire __A08_NET_194;
    wire __A08_NET_195;
    wire __A08_NET_196;
    wire __A08_NET_197;
    wire __A08_NET_198;
    wire __A08_NET_199;
    wire __A08_NET_200;
    wire __A08_NET_205;
    wire __A08_NET_206;
    wire __A08_NET_207;
    wire __A08_NET_209;
    wire __A08_NET_210;
    wire __A08_NET_211;
    wire __A08_NET_212;
    wire __A08_NET_213;
    wire __A08_NET_214;
    wire __A08_NET_215;
    wire __A08_NET_216;
    wire __A08_NET_219;
    wire __A08_NET_220;
    wire __A08_NET_221;
    wire __A08_NET_222;
    wire __A08_NET_223;
    wire __A08_NET_224;
    wire __A08_NET_225;
    wire __A08_NET_226;
    wire __A08_NET_227;
    wire __A08_NET_228;
    wire __A08_NET_229;
    wire __A08_NET_230;
    wire __A08_NET_231;
    wire __A08_NET_232;
    wire __A08_NET_233;
    wire __A08_NET_234;
    wire __A08_NET_235;
    wire __A08_NET_236;
    wire __A08_NET_237;
    wire __A08_NET_238;
    wire __A08_NET_239;
    wire __A08_NET_240;
    wire __A08_NET_241;
    wire __A08_NET_242;
    wire __A08_NET_245;
    wire __A08_NET_248;
    wire __A08_NET_249;
    wire __A08_NET_250;
    wire __A08_NET_251;
    wire __A08_NET_252;
    wire __A08_NET_253;
    wire __A08_NET_254;
    wire __A08_NET_255;
    wire __A08_NET_256;
    wire __A08_NET_257;
    wire __A08_NET_260;
    wire __A08_NET_261;
    wire __A08_NET_262;
    wire __A08_NET_263;
    wire __A08_NET_268;
    wire __A08_NET_269;
    wire __A08_NET_270;
    wire __A08_NET_271;
    wire __A08_NET_272;
    wire __A08_NET_273;
    wire __A08_NET_274;
    wire __A08_NET_275;
    wire __A08_NET_276;
    wire __A08_NET_277;
    wire __A08_NET_278;
    wire __A08_NET_279;
    wire __A08_NET_280;
    wire __A08_NET_281;
    wire __A08_NET_282;
    wire __A08_NET_283;
    wire __A08_NET_284;
    wire __A08_NET_285;
    wire __A08_NET_286;
    wire __A08_NET_287;
    wire __A08_NET_288;
    wire __A08_NET_289;
    wire __A08_NET_290;
    wire __A08_NET_291;
    wire __A08_NET_293;
    wire __A08_NET_294;
    wire __A08_NET_298;
    wire __A08_NET_299;
    wire __A08_NET_300;
    wire __A08_NET_302;
    wire __A08_NET_303;
    wire __A08_NET_304;
    wire __A08_NET_305;
    wire __A08_NET_306;
    wire __A08_NET_307;
    wire __A08_NET_308;
    wire __A08_NET_309;
    wire __A08_NET_312;
    wire __A08_NET_313;
    wire __A08_NET_314;
    wire __A08_NET_315;
    wire __A08_NET_316;
    wire __A08_NET_317;
    wire __A08_NET_318;
    wire __A08_NET_319;
    wire __A08_NET_320;
    wire __A08_NET_321;
    wire __A08_NET_322;

    pullup R8001(__A08_2___CO_IN);
    pullup R8002(RL01_n);
    pullup R8003(L01_n);
    pullup R8005(__A08_1___Z1_n);
    pullup R8006(G01_n);
    pullup R8007(RL02_n);
    pullup R8008(L02_n);
    pullup R8009(__A08_1___Z2_n);
    pullup R8010(__A08_1___G2_n);
    pullup R8011(CO06);
    pullup R8012(RL03_n);
    pullup R8013(__A08_2___L1_n);
    pullup R8015(__A08_2___Z1_n);
    pullup R8016(__A08_2___G1_n);
    pullup R8017(RL04_n);
    pullup R8018(L04_n);
    pullup R8019(__A08_2___Z2_n);
    pullup R8020(__A08_2___G2_n);
    U74HC02 U8001(__A08_NET_205, A2XG_n, __A08_1___A1_n, __A08_NET_200, WYLOG_n, WL01_n, GND, WL16_n, WYDLOG_n, __A08_NET_199, __A08_1__Y1_n, CUG, __A08_1__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8002(PONEX, __A08_NET_205, __A08_1__X1_n, CLXC, CUG, __A08_1__X1, GND, __A08_1__Y1_n, __A08_NET_200, __A08_NET_199, __A08_1__Y1, __A08_1__X1_n, __A08_1__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8003(__A08_NET_209, __A08_1__X1_n, __A08_1__Y1_n, XUY01_n, __A08_1__X1, __A08_1__Y1, GND, __A08_NET_209, XUY01_n, __A08_NET_207, __A08_NET_209, SUMA01_n, __A08_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8004( ,  , SUMA01_n, SUMB01_n, RULOG_n, __A08_NET_187, GND, __A08_NET_191, __A08_2___XUY1, XUY01_n, CI01_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U8005(CI01_n, __A08_NET_206, G01_n, GEM01, RL01_n, WL01, GND, WL01_n, WL01, __A08_1___MWL1, RL01_n, __A08_NET_157, __A08_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8006(SUMB01_n, __A08_NET_207, __A08_NET_206, __A08_NET_190, WAG_n, WL01_n, GND, WL03_n, WALSG_n, __A08_NET_192, __A08_1___A1_n, CAG, __A08_NET_188, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U8007(__A08_NET_191, __A08_2___CO_IN, __A08_NET_185, RL01_n, __A08_NET_198, L01_n, GND, __A08_1___Z1_n, __A08_NET_221, RL01_n, __A08_NET_222, RL01_n, __A08_NET_220, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U8008(__A08_NET_186, RAG_n, __A08_1___A1_n, __A08_NET_189, WLG_n, WL01_n, GND, __A08_2___G2_n, G2LSG_n, __A08_NET_196, L01_n, CLG1G, __A08_NET_197, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8009( ,  ,  , __A08_NET_194, WQG_n, WL01_n, GND, __A08_NET_194, __A08_NET_193, __A08_1___Q1_n, __A08_1___Q1_n, CQG, __A08_NET_193, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8010(__A08_NET_195, RQG_n, __A08_1___Q1_n, __A08_NET_224, WZG_n, WL01_n, GND, __A08_NET_224, __A08_NET_223, __A08_NET_221, __A08_1___Z1_n, CZG, __A08_NET_223, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8011(__A08_1___RL_OUT_1, __A08_NET_195, MDT01, RB1, R15, __A08_NET_220, GND, __A08_NET_227, __A08_NET_225, __A08_NET_226, __A08_NET_212, __A08_NET_222, __A08_NET_219, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8012(__A08_NET_219, RZG_n, __A08_1___Z1_n, __A08_NET_228, WBG_n, WL01_n, GND, __A08_NET_228, __A08_NET_229, __A08_1___B1_n, __A08_1___B1_n, CBG, __A08_NET_229, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U8013(__A08_NET_170, __A08_2___CO_IN, __A08_NET_227, RL01_n, __A08_NET_211, G01_n, GND, G01_n, __A08_NET_210, RL02_n, __A08_NET_137, L02_n, __A08_NET_147, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U8014(__A08_NET_225, RBLG_n, __A08_1___B1_n, __A08_NET_226, __A08_NET_229, RCG_n, GND, WL16_n, WG3G_n, __A08_NET_216, WL02_n, WG4G_n, __A08_NET_215, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8015(__A08_NET_190, __A08_NET_192, __A08_NET_187, __A08_NET_186, CH01, __A08_NET_185, GND, __A08_NET_198, __A08_NET_189, __A08_NET_196, __A08_NET_197, __A08_1___A1_n, __A08_NET_188, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8016(__A08_NET_214, L2GDG_n, MCRO_n, __A08_NET_213, WG1G_n, WL01_n, GND, G01_n, CGG, G01, RGG_n, G01_n, __A08_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U8017(__A08_NET_214, __A08_NET_213, WHOMPA, __A08_2___XUY2, XUY02_n, __A08_NET_170, GND, __A08_1___RL_OUT_1, RLG_n, L01_n, GND, __A08_NET_210, G01, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U8018(__A08_NET_211, G01ED, SA01, __A08_NET_216, __A08_NET_215,  , GND,  , G02ED, SA02, __A08_NET_164, __A08_NET_163, __A08_NET_162, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8019(__A08_NET_158, A2XG_n, __A08_1___A2_n, __A08_NET_160, WYLOG_n, WL02_n, GND, WL01_n, WYDG_n, __A08_NET_159, __A08_1__Y2_n, CUG, __A08_1__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8020(TWOX, __A08_NET_158, __A08_1__X2_n, CLXC, CUG, __A08_1__X2, GND, __A08_1__Y2_n, __A08_NET_160, __A08_NET_159, __A08_1__Y2, __A08_1__X2_n, __A08_1__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8021(__A08_NET_152, __A08_1__X2_n, __A08_1__Y2_n, XUY02_n, __A08_1__X2, __A08_1__Y2, GND,  ,  ,  , __A08_NET_152, XUY02_n, __A08_NET_155, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8022( ,  , __A08_NET_152, SUMA02_n, GND, __A08_2___CI_IN, GND, __A08_NET_156, SUMA02_n, SUMB02_n, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U8023(SUMB02_n, __A08_NET_155, __A08_NET_157, __A08_NET_141, WAG_n, WL02_n, GND, WL04_n, WALSG_n, __A08_NET_140, __A08_1___A2_n, CAG, __A08_NET_139, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8024(__A08_NET_141, __A08_NET_140, __A08_NET_156, __A08_NET_142, CH02, __A08_NET_137, GND, __A08_NET_147, __A08_NET_175, __A08_NET_176, __A08_NET_177, __A08_1___A2_n, __A08_NET_139, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8025(__A08_NET_142, RAG_n, __A08_1___A2_n, __A08_NET_175, WLG_n, WL02_n, GND, G05_n, G2LSG_n, __A08_NET_176, L02_n, CLG1G, __A08_NET_177, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8026(RLG_n, L02_n, __A08_1___RL_OUT_2, __A08_NET_143, __A08_NET_149, __A08_NET_148, GND, __A08_NET_138, MDT02, R1C, RB2, __A08_1___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8027(__A08_NET_179, WQG_n, WL02_n, __A08_1___Q2_n, __A08_NET_179, __A08_NET_178, GND, __A08_1___Q2_n, CQG, __A08_NET_178, RQG_n, __A08_1___Q2_n, __A08_NET_143, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U8028(__A08_NET_148, RL02_n, __A08_NET_145, __A08_1___Z2_n, __A08_NET_138, RL02_n, GND, RL02_n, __A08_NET_180, __A08_1___G2_n, __A08_NET_162, __A08_1___G2_n, __A08_NET_169, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8029(__A08_NET_144, WZG_n, WL02_n, __A08_NET_145, __A08_NET_144, __A08_NET_146, GND, __A08_1___Z2_n, CZG, __A08_NET_146, RZG_n, __A08_1___Z2_n, __A08_NET_149, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8030(__A08_NET_183, WBG_n, WL02_n, __A08_1___B2_n, __A08_NET_183, __A08_NET_184, GND, __A08_1___B2_n, CBG, __A08_NET_184, RBLG_n, __A08_1___B2_n, __A08_NET_182, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U8031(__A08_NET_182, __A08_NET_181, __A08_NET_168, __A08_NET_167, G02, __A08_NET_169, GND, __A08_NET_263, GND, XUY06_n, __A08_2___XUY2, __A08_NET_180, __A08_NET_161, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8032(__A08_NET_181, __A08_NET_184, RCG_n, __A08_NET_164, WL01_n, WG3G_n, GND, WL03_n, WG4G_n, __A08_NET_163, L2GDG_n, L01_n, __A08_NET_168, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8033(__A08_NET_167, WG1G_n, WL02_n, G02, __A08_1___G2_n, CGG, GND, RGG_n, __A08_1___G2_n, __A08_NET_161,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U8034(__A08_1___G2_n, GEM02, RL02_n, WL02, WL02, WL02_n, GND, __A08_1___MWL2, RL02_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U8035(__A08_NET_298, A2XG_n, __A08_2___A1_n, __A08_NET_294, WYLOG_n, WL03_n, GND, WL02_n, WYDG_n, __A08_NET_293, __A08_2__Y1_n, CUG, __A08_2__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8036(MONEX, __A08_NET_298, __A08_2__X1_n, CLXC, CUG, __A08_2__X1, GND, __A08_2__Y1_n, __A08_NET_294, __A08_NET_293, __A08_2__Y1, __A08_2__X1_n, __A08_2__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8037(__A08_NET_302, __A08_2__X1_n, __A08_2__Y1_n, __A08_2___XUY1, __A08_2__X1, __A08_2__Y1, GND, __A08_NET_302, __A08_2___XUY1, __A08_NET_299, __A08_NET_302, SUMA03_n, __A08_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8038( ,  , SUMA03_n, SUMB03_n, RULOG_n, __A08_NET_280, GND, __A08_NET_284, XUY05_n, __A08_2___XUY1, __A08_2___CI_IN,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U8039(__A08_2___CI_IN, __A08_NET_300, __A08_2___G1_n, GEM03, RL03_n, WL03, GND, WL03_n, WL03, __A08_2___MWL1, RL03_n, __A08_NET_250, __A08_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8040(SUMB03_n, __A08_NET_299, __A08_NET_300, __A08_NET_283, WAG_n, WL03_n, GND, WL05_n, WALSG_n, __A08_NET_285, __A08_2___A1_n, CAG, __A08_NET_281, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U8041(__A08_NET_284, CO06, __A08_NET_279, RL03_n, __A08_NET_291, __A08_2___L1_n, GND, __A08_2___Z1_n, __A08_NET_314, RL03_n, __A08_NET_315, RL03_n, __A08_NET_313, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 #(1'b1, 1'b0, 1'b1) U8042(__A08_NET_283, __A08_NET_285, __A08_NET_280, __A08_NET_278, CH03, __A08_NET_279, GND, __A08_NET_291, __A08_NET_282, __A08_NET_289, __A08_NET_290, __A08_2___A1_n, __A08_NET_281, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8043(__A08_NET_278, RAG_n, __A08_2___A1_n, __A08_NET_282, WLG_n, WL03_n, GND, G06_n, G2LSG_n, __A08_NET_289, __A08_2___L1_n, CLG1G, __A08_NET_290, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8044( ,  ,  ,  ,  ,  , GND, __A08_2___RL_OUT_1, RLG_n, __A08_2___L1_n, GND,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8045( ,  ,  , __A08_NET_287, WQG_n, WL03_n, GND, __A08_NET_287, __A08_NET_286, __A08_2___Q1_n, __A08_2___Q1_n, CQG, __A08_NET_286, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8046(__A08_NET_288, RQG_n, __A08_2___Q1_n, __A08_NET_317, WZG_n, WL03_n, GND, __A08_NET_317, __A08_NET_316, __A08_NET_314, __A08_2___Z1_n, CZG, __A08_NET_316, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8047(__A08_NET_312, RZG_n, __A08_2___Z1_n, __A08_NET_321, WBG_n, WL03_n, GND, __A08_NET_321, __A08_NET_322, __A08_2___B1_n, __A08_2___B1_n, CBG, __A08_NET_322, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8048(__A08_NET_319, RBLG_n, __A08_2___B1_n, __A08_NET_320, __A08_NET_322, RCG_n, GND, WL02_n, WG3G_n, __A08_NET_309, WL04_n, WG4G_n, __A08_NET_308, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8049(__A08_2___RL_OUT_1, __A08_NET_288, MDT03, R1C, R15, __A08_NET_313, GND, __A08_NET_318, __A08_NET_319, __A08_NET_320, __A08_NET_305, __A08_NET_315, __A08_NET_312, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U8050(__A08_NET_263, CO06, __A08_NET_318, RL03_n, __A08_NET_304, __A08_2___G1_n, GND, __A08_2___G1_n, __A08_NET_303, RL04_n, __A08_NET_230, L04_n, __A08_NET_240, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 U8051(__A08_NET_307, L2GDG_n, L02_n, __A08_NET_306, WG1G_n, WL03_n, GND, __A08_2___G1_n, CGG, G03, RGG_n, __A08_2___G1_n, __A08_NET_305, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U8052(__A08_NET_304, G03ED, SA03, __A08_NET_309, __A08_NET_308,  , GND,  , G04ED, SA04, __A08_NET_257, __A08_NET_256, __A08_NET_255, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U8053(__A08_NET_307, __A08_NET_306,  ,  ,  ,  , GND,  ,  ,  ,  , __A08_NET_303, G03, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8054(__A08_NET_251, A2XG_n, __A08_2___A2_n, __A08_NET_253, WYLOG_n, WL04_n, GND, WL03_n, WYDG_n, __A08_NET_252, __A08_2__Y2_n, CUG, __A08_2__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8055(MONEX, __A08_NET_251, __A08_2__X2_n, CLXC, CUG, __A08_2__X2, GND, __A08_2__Y2_n, __A08_NET_253, __A08_NET_252, __A08_2__Y2, __A08_2__X2_n, __A08_2__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8056(__A08_NET_245, __A08_2__X2_n, __A08_2__Y2_n, __A08_2___XUY2, __A08_2__X2, __A08_2__Y2, GND,  ,  ,  , __A08_NET_245, __A08_2___XUY2, __A08_NET_248, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8057( ,  , __A08_NET_245, __A08_2___SUMA2, __A08_2___CO_IN, CI05_n, GND, __A08_NET_249, __A08_2___SUMA2, __A08_2___SUMB2, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U8058(__A08_2___SUMB2, __A08_NET_248, __A08_NET_250, __A08_NET_234, WAG_n, WL04_n, GND, WL06_n, WALSG_n, __A08_NET_233, __A08_2___A2_n, CAG, __A08_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8059(__A08_NET_234, __A08_NET_233, __A08_NET_249, __A08_NET_235, CH04, __A08_NET_230, GND, __A08_NET_240, __A08_NET_268, __A08_NET_269, __A08_NET_270, __A08_2___A2_n, __A08_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8060(__A08_NET_235, RAG_n, __A08_2___A2_n, __A08_NET_268, WLG_n, WL04_n, GND, G07_n, G2LSG_n, __A08_NET_269, L04_n, CLG1G, __A08_NET_270, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8061(RLG_n, L04_n, __A08_2___RL_OUT_2, __A08_NET_236, __A08_NET_242, __A08_NET_241, GND, __A08_NET_231, MDT04, R1C, R15, __A08_2___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8062(__A08_NET_272, WQG_n, WL04_n, __A08_2___Q2_n, __A08_NET_272, __A08_NET_271, GND, __A08_2___Q2_n, CQG, __A08_NET_271, RQG_n, __A08_2___Q2_n, __A08_NET_236, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U8063(__A08_NET_241, RL04_n, __A08_NET_238, __A08_2___Z2_n, __A08_NET_231, RL04_n, GND, RL04_n, __A08_NET_273, __A08_2___G2_n, __A08_NET_255, __A08_2___G2_n, __A08_NET_262, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8064(__A08_NET_237, WZG_n, WL04_n, __A08_NET_238, __A08_NET_237, __A08_NET_239, GND, __A08_2___Z2_n, CZG, __A08_NET_239, RZG_n, __A08_2___Z2_n, __A08_NET_242, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8065(__A08_NET_276, WBG_n, WL04_n, __A08_2___B2_n, __A08_NET_276, __A08_NET_277, GND, __A08_2___B2_n, CBG, __A08_NET_277, RBLG_n, __A08_2___B2_n, __A08_NET_275, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U8066(__A08_NET_275, __A08_NET_274, __A08_NET_261, __A08_NET_260, G04, __A08_NET_262, GND,  ,  ,  ,  , __A08_NET_273, __A08_NET_254, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8067(__A08_NET_274, __A08_NET_277, RCG_n, __A08_NET_257, WL03_n, WG3G_n, GND, WL05_n, WG4G_n, __A08_NET_256, L2GDG_n, __A08_2___L1_n, __A08_NET_261, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8068(__A08_NET_260, WG1G_n, WL04_n, G04, __A08_2___G2_n, CGG, GND, RGG_n, __A08_2___G2_n, __A08_NET_254,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U8069(__A08_2___G2_n, GEM04, RL04_n, WL04, WL04, WL04_n, GND, __A08_2___MWL2, RL04_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC4002 U8070(SUMA01_n, __A08_NET_209, XUY01_n, CI01_n, GND,  , GND,  , __A08_NET_152, XUY02_n, __A08_1___CI_INTERNAL, WHOMP, SUMA02_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U8071(SUMA03_n, __A08_NET_302, __A08_2___XUY1, __A08_2___CI_IN, GND,  , GND,  , __A08_NET_245, __A08_2___XUY2, __A08_2___CI_INTERNAL, WHOMP, __A08_2___SUMA2, VCC, SIM_RST, SIM_CLK);
endmodule