`timescale 1ns/1ps

module agc(VCC, GND, SIM_RST, ALGA, C24A, C25A, C26A, C27A, C30A, C37P, C40P, C41P, C42P, C43P, C44P, CDUSTB_n, CHINC_n, CLOCK, CYL_n, CYR_n, DINC, DINC_n, EAC_n, EDOP_n, EXTPLS, FETCH0, FETCH0_n, FETCH1, GEQZRO_n, GINH, INCSET_n, INHPLS, INKL, INKL_n, INOTLD, L01_n, L02A_n, L15A_n, L15_n, MCDU, MINC, MNHRPT, MONPCH, MONWBK, MON_n, MSTP, MSTRTP, MTCSAI, OVNHRP, PCDU, PIPPLS_n, RADRG, RADRZ, RCHAT_n, RCHBT_n, RELPLS, RUPTOR_n, S11, S12, SBY, SHANC_n, SHIFT, SHIFT_n, SR_n, STBE, STBF, STFET1_n, STORE1_n, STRT1, STRT2, SUMA16_n, SUMB16_n, WL01_n, WL02_n, WL03_n, WL04_n, WL05_n, WL06_n, WL07_n, WL08_n, WL09_n, WL10_n, WL11_n, WL12_n, WL13_n, WL14_n, WL15, WL15_n, WL16, WL16_n, XB0_n, XB1_n, XB2_n, XB3_n, XB4_n, XB5_n, XB6_n, XB7_n, XT0_n, XT1_n, XT2_n, XT3_n, XT4_n, XT5_n, XT6_n, YB0_n, YT0_n);

    input wire VCC;
    input wire GND;
    input wire SIM_RST;
    input wire ALGA;
    input wire C24A;
    input wire C25A;
    input wire C26A;
    input wire C27A;
    input wire C30A;
    input wire C37P;
    input wire C40P;
    input wire C41P;
    input wire C42P;
    input wire C43P;
    input wire C44P;
    input wire CDUSTB_n;
    input wire CHINC_n;
    input wire CLOCK;
    input wire CYL_n;
    input wire CYR_n;
    input wire DINC;
    input wire DINC_n;
    input wire EAC_n;
    input wire EDOP_n;
    input wire EXTPLS;
    input wire FETCH0;
    input wire FETCH0_n;
    input wire FETCH1;
    input wire GEQZRO_n;
    input wire GINH;
    input wire INCSET_n;
    input wire INHPLS;
    input wire INKL;
    input wire INKL_n;
    input wire INOTLD;
    input wire L01_n;
    input wire L02A_n;
    input wire L15A_n;
    input wire L15_n;
    input wire MCDU;
    input wire MINC;
    input wire MNHRPT;
    input wire MONPCH;
    input wire MONWBK;
    input wire MON_n;
    input wire MSTP;
    input wire MSTRTP;
    input wire MTCSAI;
    input wire OVNHRP;
    input wire PCDU;
    input wire PIPPLS_n;
    input wire RADRG;
    input wire RADRZ;
    input wire RCHAT_n;
    input wire RCHBT_n;
    input wire RELPLS;
    input wire RUPTOR_n;
    input wire S11;
    input wire S12;
    input wire SBY;
    input wire SHANC_n;
    input wire SHIFT;
    input wire SHIFT_n;
    input wire SR_n;
    input wire STBE;
    input wire STBF;
    input wire STFET1_n;
    input wire STORE1_n;
    input wire STRT1;
    input wire STRT2;
    input wire SUMA16_n;
    input wire SUMB16_n;
    input wire WL01_n;
    input wire WL02_n;
    input wire WL03_n;
    input wire WL04_n;
    input wire WL05_n;
    input wire WL06_n;
    input wire WL07_n;
    input wire WL08_n;
    input wire WL09_n;
    input wire WL10_n;
    input wire WL11_n;
    input wire WL12_n;
    input wire WL13_n;
    input wire WL14_n;
    input wire WL15;
    input wire WL15_n;
    input wire WL16;
    input wire WL16_n;
    input wire XB0_n;
    input wire XB1_n;
    input wire XB2_n;
    input wire XB3_n;
    input wire XB4_n;
    input wire XB5_n;
    input wire XB6_n;
    input wire XB7_n;
    input wire XT0_n;
    input wire XT1_n;
    input wire XT2_n;
    input wire XT3_n;
    input wire XT4_n;
    input wire XT5_n;
    input wire XT6_n;
    input wire YB0_n;
    input wire YT0_n;
    wire CLK;
    wire CT;
    wire GOJAM_n;
    wire MGOJAM;
    wire MONEX_n;
    wire MONWT;
    wire MSTPIT_n;
    wire P01;
    wire P01_n;
    wire P02;
    wire P02_n;
    wire P03;
    wire P03_n;
    wire P04;
    wire P05;
    wire P05_n;
    wire PHS2;
    wire Q2A;
    wire RPTSET;
    wire RT;
    wire ST2_n;
    wire ST4_n;
    wire STOP;
    wire STOPA;
    wire STOP_n;
    wire TMZ_n;
    wire TSGN_n;
    wire WT;
    wire n10XP6;
    wire n5XP9;
    wire n8PP4;
    wire A2X_n;
    wire AD0;
    wire ADS0;
    wire AUG0_n;
    wire B15X;
    wire BR1;
    wire BR12B_n;
    wire BR1B2B;
    wire BR1B2B_n;
    wire BR1B2_n;
    wire BR1_n;
    wire BR2;
    wire BR2_n;
    wire BRDIF_n;
    wire CCS0;
    wire CCS0_n;
    wire CGMC;
    wire CI_n;
    wire CT_n;
    wire DAS0;
    wire DAS0_n;
    wire DAS1;
    wire DAS1_n;
    wire DCA0;
    wire DCS0;
    wire DIM0_n;
    wire DIVSTG;
    wire DIV_n;
    wire DV1;
    wire DV1376;
    wire DV1376_n;
    wire DV1_n;
    wire DV376_n;
    wire DV4;
    wire DV4B1B;
    wire DV4_n;
    wire DVST;
    wire DXCH0;
    wire EXST0_n;
    wire EXST1_n;
    wire EXT;
    wire FS01_n;
    wire GOJ1;
    wire GOJ1_n;
    wire GOJAM;
    wire IC1;
    wire IC10;
    wire IC10_n;
    wire IC11;
    wire IC11_n;
    wire IC12;
    wire IC12_n;
    wire IC13;
    wire IC14;
    wire IC15;
    wire IC15_n;
    wire IC16;
    wire IC16_n;
    wire IC17;
    wire IC2;
    wire IC2_n;
    wire IC3;
    wire IC4;
    wire IC5;
    wire IC5_n;
    wire IC6;
    wire IC7;
    wire IC8_n;
    wire IC9;
    wire INCR0;
    wire INOUT;
    wire INOUT_n;
    wire KRPT;
    wire L2GD_n;
    wire MASK0;
    wire MASK0_n;
    wire MP0;
    wire MP0T10;
    wire MP0_n;
    wire MP1;
    wire MP1_n;
    wire MP3;
    wire MP3A;
    wire MP3_n;
    wire MSU0;
    wire MSU0_n;
    wire NDR100_n;
    wire NDX0_n;
    wire NDXX1_n;
    wire NEAC;
    wire NISQ;
    wire OVF_n;
    wire P04_n;
    wire PHS2_n;
    wire PHS3_n;
    wire PHS4;
    wire PHS4_n;
    wire PIFL_n;
    wire PINC;
    wire PRINC;
    wire PTWOX;
    wire QC0_n;
    wire QC1_n;
    wire QC2_n;
    wire QC3_n;
    wire QXCH0_n;
    wire R15;
    wire R6;
    wire RAND0;
    wire RA_n;
    wire RBSQ;
    wire RB_n;
    wire RCH_n;
    wire RC_n;
    wire READ0;
    wire RG_n;
    wire RL10BB;
    wire RL_n;
    wire ROR0;
    wire RQ_n;
    wire RRPA;
    wire RSC_n;
    wire RSM3;
    wire RSM3_n;
    wire RSTSTG;
    wire RT_n;
    wire RUPT0;
    wire RUPT1;
    wire RUS_n;
    wire RU_n;
    wire RXOR0;
    wire RXOR0_n;
    wire RZ_n;
    wire SB2_n;
    wire SCAD_n;
    wire SQ0_n;
    wire SQ1_n;
    wire SQ2_n;
    wire SQEXT_n;
    wire SQR10;
    wire SQR10_n;
    wire SQR12_n;
    wire ST0_n;
    wire ST1;
    wire ST1_n;
    wire ST2;
    wire ST3_n;
    wire STD2;
    wire STRTFC;
    wire SU0;
    wire T01;
    wire T01_n;
    wire T02;
    wire T02_n;
    wire T03;
    wire T03_n;
    wire T04;
    wire T04_n;
    wire T05;
    wire T05_n;
    wire T06;
    wire T06_n;
    wire T07;
    wire T07_n;
    wire T08;
    wire T08_n;
    wire T09;
    wire T09_n;
    wire T10;
    wire T10_n;
    wire T11;
    wire T11_n;
    wire T12;
    wire T12USE_n;
    wire T12_n;
    wire TC0;
    wire TC0_n;
    wire TCF0;
    wire TCSAJ3_n;
    wire TL15;
    wire TOV_n;
    wire TPZG_n;
    wire TRSM;
    wire TS0;
    wire TS0_n;
    wire TSGU_n;
    wire TT_n;
    wire U2BBK;
    wire UNF_n;
    wire WAND0;
    wire WA_n;
    wire WB_n;
    wire WCH_n;
    wire WG_n;
    wire WL_n;
    wire WOR0;
    wire WQ_n;
    wire WSC_n;
    wire WS_n;
    wire WT_n;
    wire WY12_n;
    wire WYD_n;
    wire WY_n;
    wire WZ_n;
    wire ZAP_n;
    wire n10XP1;
    wire n10XP8;
    wire n11XP2;
    wire n1XP10;
    wire n2XP3;
    wire n2XP5;
    wire n2XP7;
    wire n2XP8;
    wire n3XP2;
    wire n3XP6;
    wire n3XP7;
    wire n4XP11;
    wire n4XP5;
    wire n5XP11;
    wire n5XP12;
    wire n5XP15;
    wire n5XP21;
    wire n5XP28;
    wire n5XP4;
    wire n6XP5;
    wire n6XP8;
    wire n7XP14;
    wire n7XP19;
    wire n7XP4;
    wire n7XP9;
    wire n8XP6;
    wire n9XP1;
    wire n9XP5;

    scaler A01(VCC, GND, SIM_RST, FS01_n, RCHAT_n, RCHBT_n);
    timer A02(VCC, GND, SIM_RST, CLOCK, MSTRTP, MSTP, PHS2, PHS2_n, PHS3_n, PHS4, PHS4_n, RT, RT_n, WT, WT_n, CT, CT_n, CLK, TT_n, P01, P01_n, P02, P02_n, P03, P03_n, P04, P04_n, P05, P05_n, SBY, ALGA, STRT1, STRT2, GOJ1, STOPA, GOJAM, GOJAM_n, STOP, STOP_n, WL15, WL15_n, WL16, WL16_n, FS01_n, T01, T01_n, T02, T02_n, T03, T03_n, T04, T04_n, T05, T05_n, T06, T06_n, T07, T07_n, T08, T08_n, T09, T09_n, T10, T10_n, T11, T11_n, T12, T12_n, OVF_n, UNF_n, SB2_n, MONWT, Q2A, MGOJAM, MSTPIT_n);
    sq_register A03(VCC, GND, SIM_RST, GOJAM, T01_n, T02, T12_n, PHS2_n, RT_n, CT_n, WT_n, WL16_n, WL14_n, WL13_n, WL12_n, WL11_n, WL10_n, INKL, INHPLS, RELPLS, OVNHRP, RUPTOR_n, RPTSET, KRPT, ST0_n, ST1_n, STD2, ST3_n, BR2_n, BR1B2B, RXOR0, EXT, EXTPLS, NISQ, n5XP4, MTCSAI, MNHRPT, RBSQ, SQ0_n, SQ1_n, SQ2_n, QC0_n, QC1_n, QC2_n, QC3_n, SQR12_n, SQR10, SQR10_n, SQEXT_n, EXST0_n, EXST1_n, STRTFC, AD0, ADS0, AUG0_n, CCS0, CCS0_n, DAS0, DAS0_n, DAS1, DAS1_n, DCA0, DCS0, DIM0_n, DXCH0, GOJ1, GOJ1_n, INCR0, MASK0, MASK0_n, MP0, MP0_n, MP1, MP1_n, MP3, MP3_n, MP3A, MSU0, MSU0_n, NDX0_n, NDXX1_n, QXCH0_n, RSM3, RSM3_n, SU0, TC0, TC0_n, TCF0, TCSAJ3_n, TS0, TS0_n, IC1, IC2, IC2_n, IC3, IC4, IC5, IC5_n, IC6, IC7, IC8_n, IC9, IC10, IC10_n, IC11, IC11_n, IC12, IC12_n, IC13, IC14, IC15, IC15_n, IC16, IC16_n, IC17);
    stage_branch A04(VCC, GND, SIM_RST, GOJAM, PHS2_n, PHS3_n, PHS4, PHS4_n, T01, T03, T01_n, T02_n, T03_n, T04_n, T05_n, T06_n, T07_n, T08_n, T09_n, T10_n, T11_n, T12_n, SQ0_n, SQ1_n, SQ2_n, QC0_n, QC1_n, QC2_n, QC3_n, SQEXT_n, SQR10, SQR10_n, SQR12_n, STRTFC, WL16_n, WL15_n, WL14_n, WL13_n, WL12_n, WL11_n, WL10_n, WL09_n, WL08_n, WL07_n, WL06_n, WL05_n, WL04_n, WL03_n, WL02_n, WL01_n, OVF_n, UNF_n, SUMA16_n, SUMB16_n, EXST0_n, EXST1_n, ST1, ST2, RSTSTG, TMZ_n, TOV_n, TSGN_n, TSGU_n, TPZG_n, DVST, GEQZRO_n, TRSM, NDR100_n, INKL, L15_n, TL15, XT1_n, XB7_n, MTCSAI, MP0_n, MP1, MP3A, MP3_n, IC12, IC13, IC15, IC15_n, TS0_n, RSM3, RSM3_n, STORE1_n, n7XP14, T12USE_n, ST0_n, ST1_n, STD2, ST3_n, ST4_n, BR1, BR1_n, BR2, BR2_n, BRDIF_n, BR12B_n, BR1B2_n, BR1B2B, BR1B2B_n, DIVSTG, KRPT, INOUT, INOUT_n, DIV_n, DV1, DV1_n, DV1376, DV1376_n, DV376_n, DV4, DV4_n, PRINC, RAND0, READ0, ROR0, RUPT0, RUPT1, RXOR0, RXOR0_n, WAND0, WOR0, B15X, CI_n, R15, RA_n, RB_n, RC_n, RSC_n, RRPA, WCH_n, WG_n, WL_n, n8PP4, n1XP10, n2XP3, n2XP5, n3XP2, n3XP7, n4XP5, n4XP11, n5XP4, n5XP11, n5XP28, n6XP5, n7XP19, n8XP6, n9XP1, MP0T10);
    crosspoint_nqi A05(VCC, GND, SIM_RST, GOJAM, T01, T01_n, T02_n, T03_n, T04_n, T05_n, T06_n, T07_n, T08_n, T09_n, T10_n, T11_n, T12, T12_n, T12USE_n, BR1, BR1_n, BR2, BR2_n, BR12B_n, BR1B2_n, BRDIF_n, S11, S12, INCSET_n, INKL_n, MONPCH, MONWBK, ADS0, CCS0, CCS0_n, CHINC_n, DAS0, DAS0_n, DAS1, DAS1_n, DV1, DV1_n, DV4, DV4_n, DIV_n, DXCH0, FETCH0, FETCH0_n, GOJ1, GOJ1_n, INOUT, INOUT_n, MASK0, MASK0_n, MP0, MP3, MP3_n, MSU0, MSU0_n, NDX0_n, PRINC, QXCH0_n, RAND0, READ0, ROR0, RSM3, RSM3_n, RUPT0, RXOR0, RXOR0_n, SHANC_n, SHIFT, SHIFT_n, STFET1_n, TC0, TC0_n, TCF0, TCSAJ3_n, TS0, TS0_n, WAND0, WOR0, IC1, IC2, IC2_n, IC3, IC4, IC5, IC5_n, IC8_n, IC9, IC10, IC10_n, IC11_n, IC12, IC12_n, IC13, IC14, IC15_n, IC16, IC16_n, C24A, C25A, C26A, C27A, C30A, C37P, C40P, C41P, C42P, C43P, C44P, XT0_n, XT2_n, XT3_n, XT4_n, XT5_n, XT6_n, YB0_n, YT0_n, n4XP5, n5XP9, n5XP11, n10XP6, A2X_n, CI_n, PINC, DVST, MONEX_n, NDR100_n, NISQ, PTWOX, R6, RA_n, RB_n, RC_n, RG_n, RL_n, RL10BB, RQ_n, RSTSTG, RU_n, RZ_n, SCAD_n, ST2_n, TMZ_n, TOV_n, TPZG_n, TSGN_n, U2BBK, WA_n, WB_n, WG_n, WL_n, WS_n, WY_n, WY12_n, WYD_n, WZ_n, DV4B1B, TRSM, n2XP7, n2XP8, n3XP6, n5XP12, n5XP15, n5XP21, n6XP8, n7XP4, n7XP9, n9XP5, n10XP1, n10XP8, n11XP2);
    crosspoint_ii A06(VCC, GND, SIM_RST, GOJAM, T01, T01_n, T02, T02_n, T03, T03_n, T04, T04_n, T05, T06, T06_n, T07, T07_n, T08, T08_n, T09, T10, T10_n, T11, T11_n, T12, T12USE_n, PHS4_n, ST2_n, BR1, BR1_n, BR2_n, BR1B2_n, BR12B_n, BR1B2B, BR1B2B_n, INKL, AD0, ADS0, AUG0_n, CCS0, CCS0_n, CDUSTB_n, DAS0, DAS1, DAS1_n, DCA0, DCS0, DIM0_n, DINC, DINC_n, DV1376, DV1376_n, DV376_n, DV4_n, DV4B1B, DXCH0, FETCH1, INCR0, INOTLD, MASK0, MCDU, MINC, MP0T10, MP1, MP1_n, MP3_n, MSU0, NDXX1_n, PCDU, PINC, PRINC, RAND0, RUPT0, RUPT1, SHIFT, STFET1_n, SU0, WAND0, IC6, IC7, IC9, IC11, IC17, B15X, DIVSTG, PTWOX, R6, R15, RADRG, RADRZ, RBSQ, RRPA, STBE, STBF, TL15, L01_n, L02A_n, L15A_n, MON_n, MONPCH, n8PP4, n1XP10, n2XP3, n2XP5, n2XP7, n2XP8, n3XP2, n3XP6, n3XP7, n4XP11, n5XP4, n5XP12, n5XP15, n5XP21, n5XP28, n6XP5, n6XP8, n7XP4, n7XP9, n7XP19, n8XP6, n9XP1, n9XP5, n10XP1, n10XP8, n11XP2, A2X_n, CGMC, CI_n, EXT, L2GD_n, MONEX_n, NEAC, PIFL_n, RB_n, RC_n, RCH_n, RG_n, RU_n, RUS_n, RZ_n, ST1, ST2, TOV_n, TSGU_n, WA_n, WB_n, WG_n, WL_n, WQ_n, WS_n, WSC_n, WY_n, WYD_n, WZ_n, ZAP_n, RPTSET, n7XP14);
    service_gates A07(VCC, GND, SIM_RST, T10_n, P04_n, CT_n, RT_n, TT_n, WT_n, MP3A, STFET1_n, A2X_n, CGMC, CI_n, L2GD_n, NEAC, PIFL_n, RA_n, RB_n, RC_n, RCH_n, RG_n, RL_n, RL10BB, RQ_n, RSC_n, RU_n, RUS_n, RZ_n, U2BBK, WA_n, WB_n, WCH_n, WG_n, WL_n, WQ_n, WS_n, WSC_n, WY_n, WY12_n, WYD_n, WZ_n, ZAP_n, CYL_n, CYR_n, EDOP_n, SR_n, EAC_n, GINH, L15_n, PIPPLS_n, SB2_n, SCAD_n, SHIFT, XB0_n, XB1_n, XB2_n, XB3_n, XB4_n, XB5_n, XB6_n, XT0_n);
endmodule
