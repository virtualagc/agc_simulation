`timescale 1ns/1ps

module crosspoint_ii(VCC, GND, SIM_RST, GOJAM, T01, T01_n, T02, T02_n, T03, T03_n, T04, T04_n, T05, T06, T06_n, T07, T07_n, T08, T08_n, T09, T10, T10_n, T11, T11_n, T12, T12USE_n, PHS4_n, ST2_n, BR1, BR1_n, BR2_n, BR1B2_n, BR12B_n, BR1B2B, BR1B2B_n, INKL, AD0, ADS0, AUG0_n, CCS0, CCS0_n, CDUSTB_n, DAS0, DAS1, DAS1_n, DCA0, DCS0, DIM0_n, DINC, DINC_n, DV1376, DV1376_n, DV376_n, DV4_n, DV4B1B, DXCH0, FETCH1, INCR0, INOTLD, MASK0, MCDU, MINC, MP0T10, MP1, MP1_n, MP3_n, MSU0, NDXX1_n, NISQ, PCDU, PINC, PRINC, RAND0, RUPT0, RUPT1, SHIFT, STFET1_n, SU0, WAND0, IC6, IC7, IC9, IC11, IC17, B15X, DIVSTG, PTWOX, R6, R15, R1C_n, RADRG, RADRZ, RB1_n, RBSQ, RRPA, STBE, STBF, TL15, L01_n, L02_n, L15_n, MON_n, MONPCH, n8PP4, n1XP10, n2XP3, n2XP5, n2XP7, n2XP8, n3XP2, n3XP6, n3XP7, n4XP11, n5XP4, n5XP12, n5XP15, n5XP21, n5XP28, n6XP5, n6XP8, n7XP4, n7XP9, n7XP19, n8XP6, n9XP1, n9XP5, n10XP1, n10XP8, n11XP2, A2X_n, BXVX, CGMC, CI_n, CLXC, EXT, L2GD_n, MCRO_n, MONEX, MONEX_n, NEAC, PIFL_n, PONEX, R1C, RB_n, RB1, RC_n, RCH_n, RG_n, RU_n, RUS_n, RZ_n, ST1, ST2, TOV_n, TSGU_n, TWOX, WA_n, WB_n, WG_n, WL_n, WQ_n, WS_n, WSC_n, WY_n, WYD_n, WZ_n, ZAP_n, RPTSET, n7XP14, WHOMP, WHOMPA);
    input wire SIM_RST;
    inout wire A2X_n;
    input wire AD0;
    input wire ADS0;
    input wire AUG0_n;
    input wire B15X;
    input wire BR1;
    input wire BR12B_n;
    input wire BR1B2B;
    input wire BR1B2B_n;
    input wire BR1B2_n;
    input wire BR1_n;
    input wire BR2_n;
    output wire BXVX;
    input wire CCS0;
    input wire CCS0_n;
    input wire CDUSTB_n;
    output wire CGMC;
    inout wire CI_n;
    output wire CLXC;
    input wire DAS0;
    input wire DAS1;
    input wire DAS1_n;
    input wire DCA0;
    input wire DCS0;
    input wire DIM0_n;
    input wire DINC;
    input wire DINC_n;
    input wire DIVSTG;
    input wire DV1376;
    input wire DV1376_n;
    input wire DV376_n;
    input wire DV4B1B;
    input wire DV4_n;
    input wire DXCH0;
    output wire EXT;
    input wire FETCH1;
    input wire GND;
    input wire GOJAM;
    input wire IC11;
    input wire IC17;
    input wire IC6;
    input wire IC7;
    input wire IC9;
    input wire INCR0;
    input wire INKL;
    input wire INOTLD;
    input wire L01_n;
    input wire L02_n;
    input wire L15_n;
    output wire L2GD_n;
    input wire MASK0;
    input wire MCDU;
    output wire MCRO_n;
    input wire MINC;
    output wire MONEX;
    inout wire MONEX_n;
    input wire MONPCH;
    input wire MON_n;
    input wire MP0T10;
    input wire MP1;
    input wire MP1_n;
    input wire MP3_n;
    input wire MSU0;
    input wire NDXX1_n;
    output wire NEAC;
    wire NET_181;
    wire NET_182;
    wire NET_184;
    wire NET_185;
    wire NET_186;
    wire NET_187;
    wire NET_188;
    wire NET_189;
    wire NET_190;
    wire NET_191;
    wire NET_192;
    wire NET_193;
    wire NET_194;
    wire NET_195;
    wire NET_196;
    wire NET_199;
    wire NET_200;
    wire NET_201;
    wire NET_202;
    wire NET_203;
    wire NET_204;
    wire NET_205;
    wire NET_206;
    wire NET_207;
    wire NET_209;
    wire NET_210;
    wire NET_211;
    wire NET_212;
    wire NET_213;
    wire NET_216;
    wire NET_217;
    wire NET_218;
    wire NET_219;
    wire NET_220;
    wire NET_221;
    wire NET_222;
    wire NET_223;
    wire NET_224;
    wire NET_225;
    wire NET_229;
    wire NET_230;
    wire NET_232;
    wire NET_233;
    wire NET_234;
    wire NET_235;
    wire NET_237;
    wire NET_239;
    wire NET_240;
    wire NET_241;
    wire NET_242;
    wire NET_243;
    wire NET_244;
    wire NET_245;
    wire NET_246;
    wire NET_247;
    wire NET_248;
    wire NET_249;
    wire NET_250;
    wire NET_251;
    wire NET_252;
    wire NET_253;
    wire NET_254;
    wire NET_256;
    wire NET_257;
    wire NET_258;
    wire NET_259;
    wire NET_260;
    wire NET_261;
    wire NET_262;
    wire NET_263;
    wire NET_264;
    wire NET_266;
    wire NET_267;
    wire NET_268;
    wire NET_269;
    wire NET_270;
    wire NET_271;
    wire NET_272;
    wire NET_273;
    wire NET_274;
    wire NET_275;
    wire NET_276;
    wire NET_277;
    wire NET_278;
    wire NET_279;
    wire NET_280;
    wire NET_281;
    wire NET_282;
    wire NET_283;
    wire NET_284;
    wire NET_285;
    wire NET_286;
    wire NET_287;
    wire NET_288;
    wire NET_289;
    wire NET_290;
    wire NET_291;
    wire NET_292;
    wire NET_293;
    wire NET_294;
    wire NET_297;
    wire NET_298;
    wire NET_299;
    wire NET_300;
    wire NET_301;
    wire NET_302;
    wire NET_303;
    wire NET_304;
    wire NET_305;
    wire NET_306;
    wire NET_307;
    wire NET_309;
    wire NET_310;
    wire NET_311;
    wire NET_312;
    wire NET_313;
    wire NET_314;
    wire NET_315;
    wire NET_316;
    wire NET_317;
    wire NET_318;
    wire NET_319;
    wire NET_320;
    wire NET_321;
    wire NET_322;
    wire NET_323;
    wire NET_324;
    wire NET_325;
    wire NET_326;
    wire NET_327;
    wire NET_328;
    wire NET_329;
    wire NET_330;
    wire NET_334;
    wire NET_335;
    wire NET_336;
    wire NET_338;
    wire NET_339;
    wire NET_340;
    wire NET_341;
    wire NET_342;
    wire NET_343;
    wire NET_344;
    wire NET_345;
    wire NET_346;
    input wire NISQ;
    input wire PCDU;
    input wire PHS4_n;
    output wire PIFL_n;
    input wire PINC;
    output wire PONEX;
    input wire PRINC;
    input wire PTWOX;
    input wire R15;
    output wire R1C;
    inout wire R1C_n;
    input wire R6;
    input wire RADRG;
    input wire RADRZ;
    input wire RAND0;
    output wire RB1;
    inout wire RB1_n;
    input wire RBSQ;
    inout wire RB_n;
    output wire RCH_n;
    inout wire RC_n;
    inout wire RG_n;
    inout wire RPTSET;
    input wire RRPA;
    input wire RUPT0;
    input wire RUPT1;
    output wire RUS_n;
    inout wire RU_n;
    inout wire RZ_n;
    input wire SHIFT;
    output wire ST1;
    output wire ST2;
    inout wire ST2_n;
    input wire STBE;
    input wire STBF;
    input wire STFET1_n;
    input wire SU0;
    input wire T01;
    input wire T01_n;
    input wire T02;
    input wire T02_n;
    input wire T03;
    input wire T03_n;
    input wire T04;
    input wire T04_n;
    input wire T05;
    input wire T06;
    input wire T06_n;
    input wire T07;
    input wire T07_n;
    input wire T08;
    input wire T08_n;
    input wire T09;
    input wire T10;
    input wire T10_n;
    input wire T11;
    input wire T11_n;
    input wire T12;
    input wire T12USE_n;
    input wire TL15;
    inout wire TOV_n;
    output wire TSGU_n;
    output wire TWOX;
    input wire VCC;
    input wire WAND0;
    inout wire WA_n;
    inout wire WB_n;
    inout wire WG_n;
    output wire WHOMP;
    output wire WHOMPA;
    inout wire WL_n;
    output wire WQ_n;
    inout wire WSC_n;
    inout wire WS_n;
    inout wire WYD_n;
    inout wire WY_n;
    inout wire WZ_n;
    output wire ZAP_n;
    wire __A06_1__DVXP1;
    wire __A06_1__L02A_n;
    wire __A06_1__L15A_n;
    wire __A06_1__RB1F;
    wire __A06_1__WHOMP_n;
    wire __A06_1__ZAP;
    wire __A06_1__ZIP;
    wire __A06_1__ZIPCI;
    wire __A06_2__10XP15;
    wire __A06_2__10XP9;
    wire __A06_2__6XP10;
    wire __A06_2__6XP12;
    wire __A06_2__7XP10;
    wire __A06_2__7XP11;
    wire __A06_2__7XP15;
    wire __A06_2__7XP7;
    wire __A06_2__8XP4;
    wire __A06_2__MOUT;
    wire __A06_2__POUT;
    wire __A06_2__PSEUDO;
    wire __A06_2__RDBANK;
    wire __A06_2__WOVR;
    wire __A06_2__ZOUT;
    input wire n10XP1;
    input wire n10XP8;
    input wire n11XP2;
    input wire n1XP10;
    input wire n2XP3;
    input wire n2XP5;
    input wire n2XP7;
    input wire n2XP8;
    input wire n3XP2;
    input wire n3XP6;
    input wire n3XP7;
    input wire n4XP11;
    input wire n5XP12;
    input wire n5XP15;
    input wire n5XP21;
    input wire n5XP28;
    input wire n5XP4;
    input wire n6XP5;
    input wire n6XP8;
    output wire n7XP14;
    input wire n7XP19;
    input wire n7XP4;
    input wire n7XP9;
    inout wire n8PP4;
    input wire n8XP6;
    input wire n9XP1;
    input wire n9XP5;

    pullup R6001(NET_287);
    pullup R6002(A2X_n);
    pullup R6003(RB_n);
    pullup R6004(WYD_n);
    pullup R6005(NET_280);
    pullup R6006(WL_n);
    pullup R6007(RG_n);
    pullup R6008(WB_n);
    pullup R6009(RU_n);
    pullup R6010(WZ_n);
    pullup R6011(TOV_n);
    pullup R6012(WSC_n);
    pullup R6013(WG_n);
    pullup R6014(NET_217);
    pullup R6015(NET_223);
    pullup R6016(MONEX_n);
    pullup R6017(RB1_n);
    pullup R6018(R1C_n);
    pullup R6019(n8PP4);
    pullup R6020(NET_203);
    pullup R6021(WS_n);
    pullup R6022(NET_206);
    pullup R6023(CI_n);
    pullup R6024(WA_n);
    pullup R6025(NET_243);
    pullup R6026(ST2_n);
    pullup R6027(RZ_n);
    pullup R6028(RC_n);
    U74HC27 U6001(T04, T07, NET_284, NET_285, NET_286, NET_283, GND, NET_301, T01, T03, T05, NET_298, T10, VCC, SIM_RST);
    U74HC02 U6002(NET_284, NET_298, DV376_n, NET_285, T01_n, DV1376_n, GND, T04_n, DV4_n, NET_286, MP1_n, NET_287, NET_288, VCC, SIM_RST);
    U74HC27 #(0, 0, 1) U6003(T07, T09, __A06_1__L15A_n, __A06_1__L02A_n, L01_n, NET_300, GND, NET_341, T05, T08, T11, NET_302, T11, VCC, SIM_RST);
    U74LVC07 U6004(NET_301, NET_287, NET_302, NET_287, NET_299, A2X_n, GND, RB_n, NET_313, WYD_n, NET_314, WY_n, NET_305, VCC, SIM_RST);
    U74HC02 #(1, 1, 1, 0) U6005(NET_312, NET_288, n2XP7, L2GD_n, __A06_1__ZIP, __A06_1__DVXP1, GND, __A06_1__DVXP1, NET_306, NET_314, NET_303, NET_304, NET_307, VCC, SIM_RST);
    U74HC04 U6006(L01_n, NET_290, __A06_1__L02A_n, NET_340, __A06_1__L15A_n, NET_289, GND, __A06_1__DVXP1, NET_283, __A06_1__ZIP, NET_312, NET_338, NET_339, VCC, SIM_RST);
    U74HC27 #(1, 0, 0) U6007(n7XP19, __A06_1__ZIP, __A06_1__DVXP1, NET_309, RBSQ, NET_313, GND, NET_316, NET_290, NET_340, NET_289, NET_299, __A06_1__DVXP1, VCC, SIM_RST);
    U74HC27 U6008(NET_289, NET_290, NET_312, NET_304, NET_303, NET_315, GND, NET_339, NET_303, NET_304, __A06_1__L02A_n, NET_304, __A06_1__L02A_n, VCC, SIM_RST);
    U74HC02 U6009(NET_306, NET_312, NET_307, NET_311, NET_312, NET_338, GND, NET_341, DV376_n, NET_310, DV1376_n, T02_n, NET_272, VCC, SIM_RST);
    U74HC04 U6010(NET_311, MCRO_n, NET_277, NET_274, NET_281, NET_282, GND, __A06_1__ZAP, ZAP_n, NET_343, NET_341, MONEX, MONEX_n, VCC, SIM_RST);
    U74HC27 U6011(NET_312, NET_338, NET_339, NET_316, NET_312, NET_309, GND, NET_303, NET_340, __A06_1__L15A_n, L01_n, __A06_1__ZIPCI, NET_300, VCC, SIM_RST);
    U74HC02 #(1, 1, 1, 0) U6012(NET_277, NET_310, NET_272, NET_281, NET_276, DIVSTG, GND, T08, T10, NET_278, MP1_n, NET_280, NET_266, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U6013(T06, T09, DV376_n, NET_275, T12USE_n, NET_276, GND, NET_279, T02, T04, T06, NET_275, T12, VCC, SIM_RST);
    U74LVC07 U6014(NET_279, NET_280, NET_278, NET_280, NET_273, WL_n, GND, RG_n, NET_270, WB_n, NET_291, RU_n, NET_292, VCC, SIM_RST);
    U74HC02 #(1, 0, 1, 0) U6015(NET_268, T01, T03, NET_267, NET_268, MP3_n, GND, NET_266, NET_267, ZAP_n, n5XP28, NET_274, TSGU_n, VCC, SIM_RST);
    U74HC02 #(1, 1, 1, 0) U6016(NET_273, NET_274, n5XP12, NET_297, RRPA, n5XP4, GND, n5XP15, n3XP6, WQ_n, n9XP5, n6XP8, NET_346, VCC, SIM_RST);
    U74HC4002 #(0, 1) U6017(NET_270, n5XP4, RADRG, NET_274, n5XP28, NET_271, GND, NET_269, n5XP28, n1XP10, NET_282, n2XP3, NET_291, VCC, SIM_RST);
    U74HC4002 U6018(NET_292, NET_282, __A06_1__ZAP, n5XP12, n6XP5, NET_293, GND, NET_294, PRINC, PINC, MINC, DINC, NET_229, VCC, SIM_RST);
    U74LVC07 U6019(NET_297, WZ_n, NET_345, TOV_n, NET_346, WSC_n, GND, WG_n, NET_342, NET_217, NET_218, NET_217, NET_219, VCC, SIM_RST);
    U74HC27 U6020(n6XP5, n3XP2, BR1_n, PHS4_n, TSGU_n, __A06_1__RB1F, GND, CLXC, TSGU_n, BR1, PHS4_n, NET_345, n9XP5, VCC, SIM_RST);
    U74HC02 #(0, 1, 1, 1) U6021(NET_342, n6XP8, n6XP8, PIFL_n, __A06_1__DVXP1, NET_344, GND, PTWOX, MONEX, NET_327, MONEX, B15X, NET_328, VCC, SIM_RST);
    U74HC27 U6022(PIFL_n, NET_343, STBE, n1XP10, STBF, NET_326, GND, NET_218, NET_263, NET_262, INCR0, NET_344, T02, VCC, SIM_RST);
    U74HC04 U6023(NET_327, TWOX, NET_328, BXVX, NET_336, NET_317, GND, NET_319, NET_317, NET_325, NET_319, NET_324, NET_325, VCC, SIM_RST);
    U74HC02 U6024(CGMC, NET_326, NET_336, NET_318, CGMC, NET_321, GND, NET_318, NET_326, NET_336, BR1, AUG0_n, NET_263, VCC, SIM_RST);
    U74HC04 #(0, 0, 0, 0, 1, 0) U6025(NET_324, NET_323, NET_323, NET_320, NET_320, NET_322, GND, NET_321, NET_322, NET_210, NET_212, NET_225, __A06_2__7XP10, VCC, SIM_RST);
    U74HC02 U6026(NET_262, DIM0_n, BR12B_n, NET_219, PINC, NET_261, GND, BR12B_n, DINC_n, NET_261, T06_n, NET_217, __A06_2__6XP10, VCC, SIM_RST);
    U74HC02 U6027(NET_222, MINC, MCDU, NET_220, AUG0_n, BR1_n, GND, DIM0_n, BR1B2B_n, NET_221, BR1B2B_n, DINC_n, NET_211, VCC, SIM_RST);
    U74HC27 U6028(NET_220, NET_221, BR1B2B_n, CDUSTB_n, DINC_n, __A06_2__POUT, GND, __A06_2__MOUT, BR12B_n, CDUSTB_n, DINC_n, NET_216, NET_211, VCC, SIM_RST);
    U74LVC07 U6029(NET_222, NET_223, NET_216, NET_223, NET_210, MONEX_n, GND, WA_n, NET_234, RB1_n, NET_225, R1C_n, NET_224, VCC, SIM_RST);
    U74HC02 U6030(NET_212, T06_n, NET_223, NET_213, PCDU, MCDU, GND, T06_n, NET_213, __A06_2__6XP12, NET_233, T07_n, NET_235, VCC, SIM_RST);
    U74HC27 #(0, 1, 1) U6031(BR2_n, DINC_n, DAS0, DAS1, MSU0, NET_233, GND, NET_234, NET_235, __A06_2__7XP7, NET_207, __A06_2__ZOUT, CDUSTB_n, VCC, SIM_RST);
    U74HC02 U6032(NET_232, DV4_n, BR1B2B, __A06_2__7XP7, T07_n, NET_237, GND, WAND0, INOTLD, NET_240, T07_n, NET_240, n7XP14, VCC, SIM_RST);
    U74HC27 U6033(NET_232, WAND0, DAS1_n, T07_n, BR1B2_n, __A06_2__7XP10, GND, __A06_2__7XP11, DAS1_n, T07_n, BR12B_n, NET_237, RAND0, VCC, SIM_RST);
    U74HC04 U6034(__A06_2__7XP11, NET_224, NET_201, PONEX, ST2_n, ST2, GND, ST1, NET_253, NET_250, __A06_2__PSEUDO, NET_251, __A06_2__RDBANK, VCC, SIM_RST);
    U74HC02 U6035(__A06_2__7XP15, NET_230, T07_n, NET_239, NET_229, T07_n, GND, PRINC, INKL, NET_186, IC9, DXCH0, NET_187, VCC, SIM_RST);
    U74HC27 U6036(PCDU, MCDU, n7XP9, n11XP2, __A06_2__7XP15, RUS_n, GND, NET_188, NET_239, NET_241, NET_207, NET_230, SHIFT, VCC, SIM_RST);
    U74LVC07 U6037(NET_188, RU_n, NET_189, WSC_n, NET_190, WG_n, GND, RB_n, NET_182, n8PP4, NET_181, n8PP4, NET_185, VCC, SIM_RST);
    U74HC27 U6038(NET_186, T07_n, T04_n, MON_n, FETCH1, NET_191, GND, NET_189, __A06_2__WOVR, NET_191, NET_192, __A06_2__WOVR, MONPCH, VCC, SIM_RST);
    U74HC02 U6039(NET_190, __A06_2__WOVR, NET_192, NET_192, T07_n, NET_187, GND, __A06_2__10XP9, NET_192, NET_182, T08_n, n8PP4, __A06_2__8XP4, VCC, SIM_RST);
    U74HC27 U6040(RUPT1, DAS1, IC17, MASK0, IC11, NET_185, GND, NET_184, IC6, IC7, IC9, NET_181, MSU0, VCC, SIM_RST);
    U74LVC07 U6041(NET_184, n8PP4, NET_204, NET_203, NET_202, NET_203, GND, WS_n, NET_205, NET_206, NET_195, NET_206, NET_194, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U6042(T08_n, RUPT0, NET_203, R6, R15, NET_205, GND, NET_194, ADS0, IC11, NET_193, NET_204, DAS0, VCC, SIM_RST);
    U74HC02 U6043(NET_202, MP1, DV1376, NET_209, MP3_n, BR1_n, GND, NET_209, CCS0, NET_195, T11_n, NET_206, NET_207, VCC, SIM_RST);
    U74HC02 U6044(NET_193, DAS1_n, BR2_n, NET_196, __A06_1__ZIPCI, __A06_2__6XP12, GND, CCS0_n, BR1B2B_n, NET_245, T10_n, NDXX1_n, EXT, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U6045(T03_n, DAS1_n, NET_248, NET_241, n2XP5, NET_260, GND, NET_257, IC7, DCS0, SU0, NET_241, ADS0, VCC, SIM_RST);
    U74HC4002 #(1, 0) U6046(NET_201, n8XP6, n7XP4, n10XP8, __A06_2__6XP10, NET_199, GND, NET_200, IC6, DCA0, AD0, NET_245, NET_246, VCC, SIM_RST);
    U74LVC07 U6047(NET_196, CI_n, NET_260, WA_n, NET_258, RC_n, GND, NET_243, NET_257, NET_243, NET_256, ST2_n, NET_259, VCC, SIM_RST);
    U74HC02 U6048(__A06_2__10XP9, T10_n, NET_246, NET_247, IC6, IC7, GND, T10_n, NET_247, NET_248, T10_n, NET_243, NET_242, VCC, SIM_RST);
    U74HC02 U6049(NET_258, NET_242, __A06_2__7XP7, NET_256, NET_244, DV4B1B, GND, CCS0_n, BR12B_n, NET_244, T10_n, MP1_n, __A06_2__10XP15, VCC, SIM_RST);
    U74HC27 U6050(__A06_2__8XP4, __A06_2__10XP15, __A06_2__8XP4, RADRZ, n9XP1, NET_252, GND, NEAC, NET_254, TL15, GOJAM, NET_259, RADRZ, VCC, SIM_RST);
    U74HC4002 U6051(NET_253, n2XP8, n10XP1, MP0T10, __A06_2__10XP15, NET_334, GND, NET_264, __A06_1__DVXP1, GOJAM, NISQ, __A06_1__WHOMP_n, WHOMP, VCC, SIM_RST);
    wire U6052_10_NC;
    wire U6052_11_NC;
    wire U6052_12_NC;
    wire U6052_13_NC;
    U74LVC07 U6052(NET_252, RZ_n, NET_250, RPTSET, NET_251, RU_n, GND, RC_n, NET_335, U6052_10_NC, U6052_11_NC, U6052_12_NC, U6052_13_NC, VCC, SIM_RST);
    U74HC02 #(1, 0, 0, 0) U6053(NET_254, MP0T10, NEAC, NET_249, RADRZ, __A06_2__PSEUDO, GND, T06_n, STFET1_n, __A06_2__RDBANK, __A06_1__ZIPCI, n3XP7, NET_335, VCC, SIM_RST);
    wire U6054_8_NC;
    wire U6054_9_NC;
    wire U6054_10_NC;
    wire U6054_11_NC;
    U74HC27 #(1, 0, 0) U6054(NET_249, GOJAM, n3XP7, n5XP21, n4XP11, RCH_n, GND, U6054_8_NC, U6054_9_NC, U6054_10_NC, U6054_11_NC, __A06_2__PSEUDO, RADRG, VCC, SIM_RST);
    U74HC04 #(0, 0, 0, 1, 0, 0) U6055(R1C_n, R1C, RB1_n, RB1, L02_n, NET_330, GND, __A06_1__L02A_n, NET_330, NET_329, L15_n, __A06_1__L15A_n, NET_329, VCC, SIM_RST);
    wire U6056_5_NC;
    wire U6056_6_NC;
    wire U6056_8_NC;
    wire U6056_9_NC;
    wire U6056_10_NC;
    wire U6056_11_NC;
    wire U6056_12_NC;
    wire U6056_13_NC;
    U74HC04 #(1, 0, 0, 0, 0, 0) U6056(NET_315, NET_305, __A06_1__WHOMP_n, WHOMPA, U6056_5_NC, U6056_6_NC, GND, U6056_8_NC, U6056_9_NC, U6056_10_NC, U6056_11_NC, U6056_12_NC, U6056_13_NC, VCC, SIM_RST);
    wire U6057_4_NC;
    wire U6057_5_NC;
    wire U6057_6_NC;
    wire U6057_8_NC;
    wire U6057_9_NC;
    wire U6057_10_NC;
    wire U6057_11_NC;
    wire U6057_12_NC;
    wire U6057_13_NC;
    U74HC02 #(1, 0, 0, 0) U6057(__A06_1__WHOMP_n, WHOMP, CLXC, U6057_4_NC, U6057_5_NC, U6057_6_NC, GND, U6057_8_NC, U6057_9_NC, U6057_10_NC, U6057_11_NC, U6057_12_NC, U6057_13_NC, VCC, SIM_RST);
endmodule