`include "components/agc_parts.v"

module sq_register(VCC, GND, SIM_RST, GOJAM, NISQ, T02, T12_n, PHS2_n, RT_n, CT_n, WT_n, WL16_n, WL14_n, WL13_n, WL12_n, WL11_n, WL10_n, EXT, EXTPLS, INKL, INKBT1, RELPLS, INHLPLS, OVNHRP, RUPTOR_n, KRPT, n5XP4, MNHRPT, MTCSAI);
    input wire SIM_RST;
    input wire CT_n;
    input wire EXT;
    input wire EXTPLS;
    input wire GND;
    input wire GOJAM;
    input wire INHLPLS;
    input wire INKBT1;
    input wire INKL;
    input wire KRPT;
    input wire MNHRPT;
    input wire MTCSAI;
    wire NET_100;
    wire NET_101;
    wire NET_102;
    wire NET_103;
    wire NET_104;
    wire NET_105;
    wire NET_106;
    wire NET_107;
    wire NET_108;
    wire NET_109;
    wire NET_110;
    wire NET_111;
    wire NET_112;
    wire NET_113;
    wire NET_114;
    wire NET_115;
    wire NET_116;
    wire NET_117;
    wire NET_118;
    wire NET_119;
    wire NET_72;
    wire NET_73;
    wire NET_74;
    wire NET_75;
    wire NET_76;
    wire NET_77;
    wire NET_78;
    wire NET_79;
    wire NET_80;
    wire NET_81;
    wire NET_82;
    wire NET_83;
    wire NET_84;
    wire NET_85;
    wire NET_86;
    wire NET_88;
    wire NET_89;
    wire NET_90;
    wire NET_91;
    wire NET_92;
    wire NET_93;
    wire NET_94;
    wire NET_95;
    wire NET_96;
    wire NET_97;
    wire NET_98;
    wire NET_99;
    input wire NISQ;
    input wire OVNHRP;
    input wire PHS2_n;
    input wire RELPLS;
    input wire RT_n;
    input wire RUPTOR_n;
    input wire T02;
    input wire T12_n;
    input wire VCC;
    input wire WL10_n;
    input wire WL11_n;
    input wire WL12_n;
    input wire WL13_n;
    input wire WL14_n;
    input wire WL16_n;
    input wire WT_n;
    wire __A03_1__CSQG;
    wire __A03_1__FUTEXT;
    wire __A03_1__IIP;
    wire __A03_1__IIP_n;
    wire __A03_1__INHINT;
    wire __A03_1__MIIP;
    wire __A03_1__MINHL;
    wire __A03_1__MSQ10;
    wire __A03_1__MSQ11;
    wire __A03_1__MSQ12;
    wire __A03_1__MSQ13;
    wire __A03_1__MSQ14;
    wire __A03_1__MSQ16;
    wire __A03_1__MSQEXT;
    wire __A03_1__NISQL;
    wire __A03_1__NISQL_n;
    wire __A03_1__QC0;
    wire __A03_1__QC0_n;
    wire __A03_1__QC1_n;
    wire __A03_1__QC2_n;
    wire __A03_1__QC3_n;
    wire __A03_1__RBSQ;
    wire __A03_1__RPTFRC;
    wire __A03_1__RPTSET;
    wire __A03_1__SQ0_n;
    wire __A03_1__SQ1_n;
    wire __A03_1__SQ2_n;
    wire __A03_1__SQ3_n;
    wire __A03_1__SQ4_n;
    wire __A03_1__SQ5;
    wire __A03_1__SQ6_n;
    wire __A03_1__SQ7_n;
    wire __A03_1__SQEXT;
    wire __A03_1__SQEXT_n;
    wire __A03_1__SQR10;
    wire __A03_1__SQR10_n;
    wire __A03_1__SQR11;
    wire __A03_1__SQR12;
    wire __A03_1__SQR12_n;
    wire __A03_1__SQR13;
    wire __A03_1__SQR14;
    wire __A03_1__SQR16;
    wire __A03_1__STRTFC;
    wire __A03_1__WSQG_n;
    wire __A03_1__wsqg;
    input wire n5XP4;

    pullup R3001(__A03_1__RPTSET);
    U74HC02 #(1, 0, 0, 0) U3001(NET_91, NISQ, __A03_1__NISQL, NET_94, __A03_1__STRTFC, NET_93, GND, RT_n, NET_88, __A03_1__RBSQ, NET_88, WT_n, __A03_1__wsqg, VCC, SIM_RST);
    U74HC27 U3002(NET_91, INKBT1, T12_n, NET_91, __A03_1__RPTFRC, NET_93, GND, __A03_1__CSQG, T12_n, CT_n, NET_94, __A03_1__NISQL, __A03_1__STRTFC, VCC, SIM_RST);
    U74HC04 U3003(__A03_1__NISQL, __A03_1__NISQL_n, NET_93, NET_88, __A03_1__wsqg, __A03_1__WSQG_n, GND, __A03_1__STRTFC, NET_86, __A03_1__SQEXT, NET_77, __A03_1__SQEXT_n, NET_76, VCC, SIM_RST);
    wire U3004_11_NC;
    wire U3004_12_NC;
    wire U3004_13_NC;
    U74HC02 U3004(NET_113, WL16_n, __A03_1__WSQG_n, NET_112, WL14_n, __A03_1__WSQG_n, GND, WL13_n, __A03_1__WSQG_n, NET_111, U3004_11_NC, U3004_12_NC, U3004_13_NC, VCC, SIM_RST);
    U74HC02 U3005(NET_86, GOJAM, MTCSAI, NET_90, __A03_1__NISQL_n, T12_n, GND, __A03_1__STRTFC, NET_90, NET_75, NET_75, NET_89, NET_74, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U3006(EXTPLS, EXT, NET_89, INKBT1, __A03_1__STRTFC, __A03_1__FUTEXT, GND, NET_77, __A03_1__RPTFRC, NET_74, NET_76, NET_89, __A03_1__FUTEXT, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 1) U3007(NET_73, NET_75, __A03_1__FUTEXT, NET_76, NET_77, NET_73, GND, INHLPLS, __A03_1__INHINT, NET_72, KRPT, __A03_1__IIP, __A03_1__IIP_n, VCC, SIM_RST);
    U74HC04 U3008(NET_77, __A03_1__MSQEXT, NET_72, __A03_1__MINHL, __A03_1__IIP_n, __A03_1__MIIP, GND, __A03_1__MSQ16, NET_102, __A03_1__MSQ14, NET_117, __A03_1__MSQ13, NET_118, VCC, SIM_RST);
    U74HC27 U3009(NET_72, RELPLS, __A03_1__IIP_n, GOJAM, n5XP4, __A03_1__IIP, GND, NET_82, __A03_1__FUTEXT, __A03_1__NISQL_n, T12_n, __A03_1__INHINT, GOJAM, VCC, SIM_RST);
    U74HC27 U3010(PHS2_n, RUPTOR_n, OVNHRP, __A03_1__INHINT, __A03_1__IIP, NET_80, GND, NET_78, NET_79, __A03_1__STRTFC, T02, NET_81, MNHRPT, VCC, SIM_RST);
    wire U3011_8_NC;
    wire U3011_9_NC;
    wire U3011_10_NC;
    wire U3011_11_NC;
    wire U3011_12_NC;
    wire U3011_13_NC;
    U74LVC07 U3011(NET_82, __A03_1__RPTSET, NET_81, __A03_1__RPTSET, NET_80, __A03_1__RPTSET, GND, U3011_8_NC, U3011_9_NC, U3011_10_NC, U3011_11_NC, U3011_12_NC, U3011_13_NC, VCC, SIM_RST);
    U74HC02 #(1, 1, 1, 1) U3012(NET_79, __A03_1__RPTSET, NET_78, NET_102, NET_113, __A03_1__SQR16, GND, NET_112, __A03_1__SQR14, NET_117, NET_111, __A03_1__SQR13, NET_118, VCC, SIM_RST);
    U74HC27 U3013(NET_102, __A03_1__RPTFRC, NET_117, __A03_1__RPTFRC, __A03_1__CSQG, __A03_1__SQR14, GND, __A03_1__SQR13, NET_118, __A03_1__RPTFRC, __A03_1__CSQG, __A03_1__SQR16, __A03_1__CSQG, VCC, SIM_RST);
    wire U3014_8_NC;
    wire U3014_9_NC;
    wire U3014_10_NC;
    wire U3014_11_NC;
    wire U3014_12_NC;
    wire U3014_13_NC;
    U74HC02 U3014(NET_101, NET_102, INKL, NET_100, INKL, __A03_1__SQR16, GND, U3014_8_NC, U3014_9_NC, U3014_10_NC, U3014_11_NC, U3014_12_NC, U3014_13_NC, VCC, SIM_RST);
    U74HC27 U3015(NET_115, NET_119, NET_118, NET_119, NET_104, NET_109, GND, NET_108, NET_115, NET_117, NET_104, NET_110, NET_104, VCC, SIM_RST);
    U74HC27 U3016(NET_118, NET_117, NET_115, NET_119, NET_114, NET_106, GND, __A03_1__SQ5, NET_118, NET_119, NET_114, NET_107, NET_104, VCC, SIM_RST);
    U74HC27 #(0, 0, 1) U3017(NET_115, NET_114, NET_118, NET_117, NET_114, NET_103, GND, NET_83, __A03_1__RPTFRC, NET_116, __A03_1__SQR12, NET_105, NET_117, VCC, SIM_RST);
    U74HC04 U3018(NET_109, __A03_1__SQ1_n, NET_108, __A03_1__SQ2_n, NET_107, __A03_1__SQ3_n, GND, __A03_1__SQ4_n, NET_106, __A03_1__SQ6_n, NET_105, __A03_1__SQ7_n, NET_103, VCC, SIM_RST);
    U74HC02 U3019(NET_116, WL12_n, __A03_1__WSQG_n, NET_85, WL11_n, __A03_1__WSQG_n, GND, NET_83, __A03_1__CSQG, __A03_1__SQR12, NET_84, __A03_1__CSQG, __A03_1__SQR11, VCC, SIM_RST);
    wire U3020_8_NC;
    wire U3020_9_NC;
    wire U3020_10_NC;
    wire U3020_11_NC;
    U74HC27 #(1, 1, 0) U3020(__A03_1__RPTFRC, NET_85, __A03_1__RPTFRC, NET_99, NET_98, NET_97, GND, U3020_8_NC, U3020_9_NC, U3020_10_NC, U3020_11_NC, NET_84, __A03_1__SQR11, VCC, SIM_RST);
    wire U3021_12_NC;
    wire U3021_13_NC;
    U74HC04 U3021(NET_83, __A03_1__MSQ12, NET_84, __A03_1__MSQ11, NET_97, __A03_1__MSQ10, GND, __A03_1__SQR12_n, __A03_1__SQR12, __A03_1__RPTFRC, NET_79, U3021_12_NC, U3021_13_NC, VCC, SIM_RST);
    U74HC02 U3022(__A03_1__QC0, __A03_1__SQR11, __A03_1__SQR12, NET_95, NET_84, __A03_1__SQR12, GND, __A03_1__SQR11, NET_83, NET_92, NET_83, NET_84, NET_96, VCC, SIM_RST);
    U74HC04 U3023(__A03_1__QC0, __A03_1__QC0_n, NET_95, __A03_1__QC1_n, NET_92, __A03_1__QC2_n, GND, __A03_1__QC3_n, NET_96, __A03_1__SQR10, NET_97, __A03_1__SQR10_n, NET_98, VCC, SIM_RST);
    wire U3024_8_NC;
    wire U3024_9_NC;
    wire U3024_10_NC;
    wire U3024_11_NC;
    wire U3024_12_NC;
    wire U3024_13_NC;
    U74HC02 U3024(NET_99, WL10_n, __A03_1__WSQG_n, NET_98, NET_97, __A03_1__CSQG, GND, U3024_8_NC, U3024_9_NC, U3024_10_NC, U3024_11_NC, U3024_12_NC, U3024_13_NC, VCC, SIM_RST);
    wire U3025_12_NC;
    wire U3025_13_NC;
    U74HC04 U3025(NET_101, NET_114, NET_100, NET_104, NET_117, NET_119, GND, NET_115, NET_118, __A03_1__SQ0_n, NET_110, U3025_12_NC, U3025_13_NC, VCC, SIM_RST);
endmodule