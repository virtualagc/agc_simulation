`timescale 1ns/1ps

module four_bit_3(VCC, GND, SIM_RST, A2XG_n, CAG, CBG, CGG, CLG1G, CLXC, CQG, CUG, CZG, L2GDG_n, RAG_n, RCG_n, RGG_n, RLG_n, RQG_n, RZG_n, WAG_n, WALSG_n, WBG_n, WLG_n, WQG_n, WZG_n, CI09_n, CO10, MONEX, XUY13_n, XUY14_n, CH09, CH10, CH11, CH12, L08_n, G2LSG_n, G13_n, G14_n, G15_n, MDT09, MDT10, MDT11, MDT12, SA09, SA10, SA11, SA12, RBHG_n, RBLG_n, RULOG_n, WL13_n, WL14_n, WG1G_n, WG3G_n, WG4G_n, WYDG_n, WYLOG_n, R1C, WL08_n, G09_n, G10_n, G11_n, WL09_n, WL10_n, WL11_n, WL12_n, XUY09_n, XUY10_n);
    input wire SIM_RST;
    input wire A2XG_n;
    input wire CAG;
    input wire CBG;
    input wire CGG;
    input wire CH09;
    input wire CH10;
    input wire CH11;
    input wire CH12;
    input wire CI09_n;
    input wire CLG1G;
    input wire CLXC;
    input wire CO10;
    input wire CQG;
    input wire CUG;
    input wire CZG;
    inout wire G09_n;
    inout wire G10_n;
    inout wire G11_n;
    input wire G13_n;
    input wire G14_n;
    input wire G15_n;
    input wire G2LSG_n;
    input wire GND;
    input wire L08_n;
    input wire L2GDG_n;
    input wire MDT09;
    input wire MDT10;
    input wire MDT11;
    input wire MDT12;
    input wire MONEX;
    wire NET_123;
    wire NET_124;
    wire NET_125;
    wire NET_126;
    wire NET_127;
    wire NET_128;
    wire NET_129;
    wire NET_130;
    wire NET_131;
    wire NET_132;
    wire NET_133;
    wire NET_136;
    wire NET_137;
    wire NET_138;
    wire NET_139;
    wire NET_140;
    wire NET_141;
    wire NET_142;
    wire NET_146;
    wire NET_147;
    wire NET_148;
    wire NET_149;
    wire NET_150;
    wire NET_151;
    wire NET_152;
    wire NET_153;
    wire NET_154;
    wire NET_157;
    wire NET_158;
    wire NET_159;
    wire NET_160;
    wire NET_161;
    wire NET_162;
    wire NET_163;
    wire NET_164;
    wire NET_165;
    wire NET_166;
    wire NET_167;
    wire NET_168;
    wire NET_169;
    wire NET_170;
    wire NET_171;
    wire NET_172;
    wire NET_173;
    wire NET_174;
    wire NET_175;
    wire NET_176;
    wire NET_177;
    wire NET_178;
    wire NET_179;
    wire NET_180;
    wire NET_181;
    wire NET_182;
    wire NET_183;
    wire NET_188;
    wire NET_189;
    wire NET_190;
    wire NET_191;
    wire NET_192;
    wire NET_193;
    wire NET_194;
    wire NET_195;
    wire NET_196;
    wire NET_197;
    wire NET_198;
    wire NET_199;
    wire NET_200;
    wire NET_201;
    wire NET_202;
    wire NET_203;
    wire NET_204;
    wire NET_205;
    wire NET_206;
    wire NET_207;
    wire NET_208;
    wire NET_209;
    wire NET_210;
    wire NET_211;
    wire NET_212;
    wire NET_213;
    wire NET_214;
    wire NET_215;
    wire NET_216;
    wire NET_217;
    wire NET_218;
    wire NET_219;
    wire NET_220;
    wire NET_221;
    wire NET_222;
    wire NET_223;
    wire NET_224;
    wire NET_227;
    wire NET_228;
    wire NET_229;
    wire NET_230;
    wire NET_231;
    wire NET_232;
    wire NET_233;
    wire NET_237;
    wire NET_238;
    wire NET_239;
    wire NET_240;
    wire NET_241;
    wire NET_242;
    wire NET_243;
    wire NET_244;
    wire NET_245;
    wire NET_248;
    wire NET_249;
    wire NET_250;
    wire NET_251;
    wire NET_252;
    wire NET_253;
    wire NET_254;
    wire NET_255;
    wire NET_256;
    wire NET_257;
    wire NET_258;
    wire NET_259;
    wire NET_260;
    wire NET_261;
    wire NET_262;
    wire NET_263;
    wire NET_264;
    wire NET_265;
    wire NET_266;
    wire NET_267;
    wire NET_268;
    wire NET_269;
    wire NET_270;
    wire NET_271;
    wire NET_272;
    wire NET_273;
    wire NET_274;
    wire NET_279;
    wire NET_280;
    wire NET_281;
    wire NET_282;
    wire NET_283;
    wire NET_284;
    wire NET_285;
    wire NET_286;
    wire NET_287;
    wire NET_288;
    wire NET_289;
    wire NET_290;
    wire NET_291;
    wire NET_292;
    wire NET_293;
    wire NET_294;
    wire NET_295;
    wire NET_296;
    wire NET_297;
    wire NET_298;
    wire NET_299;
    wire NET_300;
    wire NET_301;
    wire NET_302;
    wire NET_303;
    wire NET_304;
    input wire R1C;
    input wire RAG_n;
    input wire RBHG_n;
    input wire RBLG_n;
    input wire RCG_n;
    input wire RGG_n;
    input wire RLG_n;
    input wire RQG_n;
    input wire RULOG_n;
    input wire RZG_n;
    input wire SA09;
    input wire SA10;
    input wire SA11;
    input wire SA12;
    input wire VCC;
    input wire WAG_n;
    input wire WALSG_n;
    input wire WBG_n;
    input wire WG1G_n;
    input wire WG3G_n;
    input wire WG4G_n;
    input wire WL08_n;
    output wire WL09_n;
    output wire WL10_n;
    output wire WL11_n;
    output wire WL12_n;
    input wire WL13_n;
    input wire WL14_n;
    input wire WLG_n;
    input wire WQG_n;
    input wire WYDG_n;
    input wire WYLOG_n;
    input wire WZG_n;
    output wire XUY09_n;
    output wire XUY10_n;
    input wire XUY13_n;
    input wire XUY14_n;
    wire __A10_1__X1;
    wire __A10_1__X1_n;
    wire __A10_1__X2;
    wire __A10_1__X2_n;
    wire __A10_1__Y1;
    wire __A10_1__Y1_n;
    wire __A10_1__Y2;
    wire __A10_1__Y2_n;
    wire __A10_1___A1_n;
    wire __A10_1___A2_n;
    wire __A10_1___B1_n;
    wire __A10_1___B2_n;
    wire __A10_1___CI_INTERNAL;
    wire __A10_1___G1;
    wire __A10_1___G2;
    wire __A10_1___GEM1;
    wire __A10_1___GEM2;
    wire __A10_1___L1_n;
    wire __A10_1___L2_n;
    wire __A10_1___MWL1;
    wire __A10_1___MWL2;
    wire __A10_1___Q1_n;
    wire __A10_1___Q2_n;
    wire __A10_1___RL1_n;
    wire __A10_1___RL2_n;
    wire __A10_1___SUMA1;
    wire __A10_1___SUMA2;
    wire __A10_1___SUMB1;
    wire __A10_1___SUMB2;
    wire __A10_1___WL1;
    wire __A10_1___WL2;
    wire __A10_1___Z1_n;
    wire __A10_1___Z2_n;
    wire __A10_2__X1;
    wire __A10_2__X1_n;
    wire __A10_2__X2;
    wire __A10_2__X2_n;
    wire __A10_2__Y1;
    wire __A10_2__Y1_n;
    wire __A10_2__Y2;
    wire __A10_2__Y2_n;
    wire __A10_2___A1_n;
    wire __A10_2___A2_n;
    wire __A10_2___B1_n;
    wire __A10_2___B2_n;
    wire __A10_2___CI_IN;
    wire __A10_2___CI_INTERNAL;
    wire __A10_2___CI_OUT;
    wire __A10_2___CO_IN;
    wire __A10_2___CO_OUT;
    wire __A10_2___G1;
    wire __A10_2___G2;
    wire __A10_2___G2_n;
    wire __A10_2___GEM1;
    wire __A10_2___GEM2;
    wire __A10_2___L1_n;
    wire __A10_2___L2_n;
    wire __A10_2___MWL1;
    wire __A10_2___MWL2;
    wire __A10_2___Q1_n;
    wire __A10_2___Q2_n;
    wire __A10_2___RL1_n;
    wire __A10_2___RL2_n;
    wire __A10_2___SUMA1;
    wire __A10_2___SUMA2;
    wire __A10_2___SUMB1;
    wire __A10_2___SUMB2;
    wire __A10_2___WL1;
    wire __A10_2___WL2;
    wire __A10_2___XUY1;
    wire __A10_2___XUY2;
    wire __A10_2___Z1_n;
    wire __A10_2___Z2_n;

    pullup R10001(__A10_2___CO_IN);
    pullup R10002(__A10_1___RL1_n);
    pullup R10003(__A10_1___L1_n);
    pullup R10005(__A10_1___Z1_n);
    pullup R10006(G09_n);
    pullup R10007(__A10_1___RL2_n);
    pullup R10008(__A10_1___L2_n);
    pullup R10009(__A10_1___Z2_n);
    pullup R10010(G10_n);
    pullup R10011(__A10_2___CO_OUT);
    pullup R10012(__A10_2___RL1_n);
    pullup R10013(__A10_2___L1_n);
    pullup R10015(__A10_2___Z1_n);
    pullup R10016(G11_n);
    pullup R10017(__A10_2___RL2_n);
    pullup R10018(__A10_2___L2_n);
    pullup R10019(__A10_2___Z2_n);
    pullup R10020(__A10_2___G2_n);
    U74HC02 U10001(NET_188, A2XG_n, __A10_1___A1_n, NET_183, WYLOG_n, WL09_n, GND, WL08_n, WYDG_n, NET_182, __A10_1__Y1_n, CUG, __A10_1__Y1, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U10002(MONEX, NET_188, __A10_1__X1_n, CLXC, CUG, __A10_1__X1, GND, __A10_1__Y1_n, NET_183, NET_182, __A10_1__Y1, __A10_1__X1_n, __A10_1__X1, VCC, SIM_RST);
    U74HC02 U10003(NET_191, __A10_1__X1_n, __A10_1__Y1_n, XUY09_n, __A10_1__X1, __A10_1__Y1, GND, NET_191, XUY09_n, NET_190, NET_191, __A10_1___SUMA1, __A10_1___CI_INTERNAL, VCC, SIM_RST);
    U74HC27 U10004(NET_191, XUY09_n, __A10_1___SUMA1, __A10_1___SUMB1, RULOG_n, NET_173, GND, NET_175, __A10_2___XUY1, XUY09_n, CI09_n, __A10_1___SUMA1, CI09_n, VCC, SIM_RST);
    U74HC04 U10005(CI09_n, NET_189, G09_n, __A10_1___GEM1, __A10_1___RL1_n, __A10_1___WL1, GND, WL09_n, __A10_1___WL1, __A10_1___MWL1, __A10_1___RL1_n, NET_136, __A10_1___CI_INTERNAL, VCC, SIM_RST);
    U74HC02 U10006(__A10_1___SUMB1, NET_190, NET_189, NET_174, WAG_n, WL09_n, GND, WL11_n, WALSG_n, NET_171, __A10_1___A1_n, CAG, NET_170, VCC, SIM_RST);
    U74LVC07 U10007(NET_175, __A10_2___CO_IN, NET_172, __A10_1___RL1_n, NET_181, __A10_1___L1_n, GND, __A10_1___Z1_n, NET_205, __A10_1___RL1_n, NET_206, __A10_1___RL1_n, NET_212, VCC, SIM_RST);
    U74HC02 U10008(NET_169, RAG_n, __A10_1___A1_n, NET_178, WLG_n, WL09_n, GND, __A10_2___G2_n, G2LSG_n, NET_180, __A10_1___L1_n, CLG1G, NET_179, VCC, SIM_RST);
    wire U10009_1_NC;
    wire U10009_2_NC;
    wire U10009_3_NC;
    U74HC02 #(0, 0, 1, 0) U10009(U10009_1_NC, U10009_2_NC, U10009_3_NC, NET_176, WQG_n, WL09_n, GND, NET_176, NET_177, __A10_1___Q1_n, __A10_1___Q1_n, CQG, NET_177, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U10010(NET_200, RQG_n, __A10_1___Q1_n, NET_208, WZG_n, WL09_n, GND, NET_208, NET_204, NET_205, __A10_1___Z1_n, CZG, NET_204, VCC, SIM_RST);
    U74HC27 U10011(NET_210, NET_200, MDT09, R1C, GND, NET_212, GND, NET_209, NET_196, NET_195, NET_201, NET_206, NET_207, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U10012(NET_207, RZG_n, __A10_1___Z1_n, NET_213, WBG_n, WL09_n, GND, NET_213, NET_211, __A10_1___B1_n, __A10_1___B1_n, CBG, NET_211, VCC, SIM_RST);
    U74LVC07 U10013(NET_138, __A10_2___CO_IN, NET_209, __A10_1___RL1_n, NET_192, G09_n, GND, G09_n, NET_193, __A10_1___RL2_n, NET_125, __A10_1___L2_n, NET_164, VCC, SIM_RST);
    U74HC02 U10014(NET_196, RBLG_n, __A10_1___B1_n, NET_195, NET_211, RCG_n, GND, WL08_n, WG3G_n, NET_199, WL10_n, WG4G_n, NET_198, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U10015(NET_174, NET_171, NET_173, NET_169, CH09, NET_172, GND, NET_181, NET_178, NET_180, NET_179, __A10_1___A1_n, NET_170, VCC, SIM_RST);
    U74HC02 U10016(NET_197, L2GDG_n, L08_n, NET_194, WG1G_n, WL09_n, GND, G09_n, CGG, __A10_1___G1, RGG_n, G09_n, NET_201, VCC, SIM_RST);
    wire U10017_3_NC;
    wire U10017_4_NC;
    wire U10017_5_NC;
    wire U10017_6_NC;
    U74HC27 #(1, 0, 0) U10017(NET_197, NET_194, U10017_3_NC, U10017_4_NC, U10017_5_NC, U10017_6_NC, GND, NET_210, RLG_n, __A10_1___L1_n, GND, NET_193, __A10_1___G1, VCC, SIM_RST);
    U74HC4002 U10018(NET_192, GND, SA09, NET_199, NET_198, NET_203, GND, NET_202, GND, SA10, NET_149, NET_148, NET_151, VCC, SIM_RST);
    U74HC02 U10019(NET_127, A2XG_n, __A10_1___A2_n, NET_141, WYLOG_n, WL10_n, GND, WL09_n, WYDG_n, NET_142, __A10_1__Y2_n, CUG, __A10_1__Y2, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U10020(MONEX, NET_127, __A10_1__X2_n, CLXC, CUG, __A10_1__X2, GND, __A10_1__Y2_n, NET_141, NET_142, __A10_1__Y2, __A10_1__X2_n, __A10_1__X2, VCC, SIM_RST);
    U74HC02 U10021(NET_139, __A10_1__X2_n, __A10_1__Y2_n, XUY10_n, __A10_1__X2, __A10_1__Y2, GND, __A10_2___XUY2, XUY10_n, NET_138, NET_139, XUY10_n, NET_137, VCC, SIM_RST);
    U74HC27 U10022(NET_139, XUY10_n, NET_139, __A10_1___SUMA2, CO10, __A10_2___CI_IN, GND, NET_140, __A10_1___SUMA2, __A10_1___SUMB2, RULOG_n, __A10_1___SUMA2, __A10_1___CI_INTERNAL, VCC, SIM_RST);
    U74HC02 U10023(__A10_1___SUMB2, NET_137, NET_136, NET_126, WAG_n, WL10_n, GND, WL12_n, WALSG_n, NET_128, __A10_1___A2_n, CAG, NET_124, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U10024(NET_126, NET_128, NET_140, NET_123, CH10, NET_125, GND, NET_164, NET_167, NET_168, NET_160, __A10_1___A2_n, NET_124, VCC, SIM_RST);
    U74HC02 U10025(NET_123, RAG_n, __A10_1___A2_n, NET_167, WLG_n, WL10_n, GND, G13_n, G2LSG_n, NET_168, __A10_1___L2_n, CLG1G, NET_160, VCC, SIM_RST);
    U74HC27 U10026(RLG_n, __A10_1___L2_n, NET_162, NET_161, NET_129, NET_130, GND, NET_133, MDT10, R1C, GND, NET_162, GND, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U10027(NET_158, WQG_n, WL10_n, __A10_1___Q2_n, NET_158, NET_159, GND, __A10_1___Q2_n, CQG, NET_159, RQG_n, __A10_1___Q2_n, NET_161, VCC, SIM_RST);
    U74LVC07 U10028(NET_130, __A10_1___RL2_n, NET_131, __A10_1___Z2_n, NET_133, __A10_1___RL2_n, GND, __A10_1___RL2_n, NET_154, G10_n, NET_151, G10_n, NET_150, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U10029(NET_163, WZG_n, WL10_n, NET_131, NET_163, NET_132, GND, __A10_1___Z2_n, CZG, NET_132, RZG_n, __A10_1___Z2_n, NET_129, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U10030(NET_165, WBG_n, WL10_n, __A10_1___B2_n, NET_165, NET_166, GND, __A10_1___B2_n, CBG, NET_166, RBLG_n, __A10_1___B2_n, NET_153, VCC, SIM_RST);
    wire U10031_8_NC;
    wire U10031_9_NC;
    wire U10031_10_NC;
    wire U10031_11_NC;
    U74HC27 #(0, 1, 0) U10031(NET_153, NET_152, NET_147, NET_146, __A10_1___G2, NET_150, GND, U10031_8_NC, U10031_9_NC, U10031_10_NC, U10031_11_NC, NET_154, NET_157, VCC, SIM_RST);
    U74HC02 U10032(NET_152, NET_166, RCG_n, NET_149, WL09_n, WG3G_n, GND, WL11_n, WG4G_n, NET_148, L2GDG_n, __A10_1___L1_n, NET_147, VCC, SIM_RST);
    wire U10033_11_NC;
    wire U10033_12_NC;
    wire U10033_13_NC;
    U74HC02 U10033(NET_146, WG1G_n, WL10_n, __A10_1___G2, G10_n, CGG, GND, RGG_n, G10_n, NET_157, U10033_11_NC, U10033_12_NC, U10033_13_NC, VCC, SIM_RST);
    wire U10034_10_NC;
    wire U10034_11_NC;
    wire U10034_12_NC;
    wire U10034_13_NC;
    U74HC04 U10034(G10_n, __A10_1___GEM2, __A10_1___RL2_n, __A10_1___WL2, __A10_1___WL2, WL10_n, GND, __A10_1___MWL2, __A10_1___RL2_n, U10034_10_NC, U10034_11_NC, U10034_12_NC, U10034_13_NC, VCC, SIM_RST);
    U74HC02 U10035(NET_279, A2XG_n, __A10_2___A1_n, NET_274, WYLOG_n, WL11_n, GND, WL10_n, WYDG_n, NET_273, __A10_2__Y1_n, CUG, __A10_2__Y1, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U10036(MONEX, NET_279, __A10_2__X1_n, CLXC, CUG, __A10_2__X1, GND, __A10_2__Y1_n, NET_274, NET_273, __A10_2__Y1, __A10_2__X1_n, __A10_2__X1, VCC, SIM_RST);
    U74HC02 U10037(NET_282, __A10_2__X1_n, __A10_2__Y1_n, __A10_2___XUY1, __A10_2__X1, __A10_2__Y1, GND, NET_282, __A10_2___XUY1, NET_281, NET_282, __A10_2___SUMA1, __A10_2___CI_INTERNAL, VCC, SIM_RST);
    U74HC27 U10038(NET_282, __A10_2___XUY1, __A10_2___SUMA1, __A10_2___SUMB1, RULOG_n, NET_264, GND, NET_266, XUY13_n, __A10_2___XUY1, __A10_2___CI_IN, __A10_2___SUMA1, __A10_2___CI_IN, VCC, SIM_RST);
    U74HC04 U10039(__A10_2___CI_IN, NET_280, G11_n, __A10_2___GEM1, __A10_2___RL1_n, __A10_2___WL1, GND, WL11_n, __A10_2___WL1, __A10_2___MWL1, __A10_2___RL1_n, NET_227, __A10_2___CI_INTERNAL, VCC, SIM_RST);
    U74HC02 U10040(__A10_2___SUMB1, NET_281, NET_280, NET_265, WAG_n, WL11_n, GND, WL13_n, WALSG_n, NET_262, __A10_2___A1_n, CAG, NET_261, VCC, SIM_RST);
    U74LVC07 U10041(NET_266, __A10_2___CO_OUT, NET_263, __A10_2___RL1_n, NET_272, __A10_2___L1_n, GND, __A10_2___Z1_n, NET_296, __A10_2___RL1_n, NET_297, __A10_2___RL1_n, NET_303, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U10042(NET_265, NET_262, NET_264, NET_260, CH11, NET_263, GND, NET_272, NET_269, NET_271, NET_270, __A10_2___A1_n, NET_261, VCC, SIM_RST);
    U74HC02 U10043(NET_260, RAG_n, __A10_2___A1_n, NET_269, WLG_n, WL11_n, GND, G14_n, G2LSG_n, NET_271, __A10_2___L1_n, CLG1G, NET_270, VCC, SIM_RST);
    wire U10044_1_NC;
    wire U10044_2_NC;
    wire U10044_3_NC;
    wire U10044_4_NC;
    wire U10044_5_NC;
    wire U10044_6_NC;
    wire U10044_12_NC;
    wire U10044_13_NC;
    U74HC27 U10044(U10044_1_NC, U10044_2_NC, U10044_3_NC, U10044_4_NC, U10044_5_NC, U10044_6_NC, GND, NET_300, RLG_n, __A10_2___L1_n, GND, U10044_12_NC, U10044_13_NC, VCC, SIM_RST);
    wire U10045_1_NC;
    wire U10045_2_NC;
    wire U10045_3_NC;
    U74HC02 #(0, 0, 1, 0) U10045(U10045_1_NC, U10045_2_NC, U10045_3_NC, NET_267, WQG_n, WL11_n, GND, NET_267, NET_268, __A10_2___Q1_n, __A10_2___Q1_n, CQG, NET_268, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U10046(NET_283, RQG_n, __A10_2___Q1_n, NET_299, WZG_n, WL11_n, GND, NET_299, NET_295, NET_296, __A10_2___Z1_n, CZG, NET_295, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U10047(NET_298, RZG_n, __A10_2___Z1_n, NET_304, WBG_n, WL11_n, GND, NET_304, NET_302, __A10_2___B1_n, __A10_2___B1_n, CBG, NET_302, VCC, SIM_RST);
    U74HC02 U10048(NET_288, RBHG_n, __A10_2___B1_n, NET_287, NET_302, RCG_n, GND, WL10_n, WG3G_n, NET_291, WL12_n, WG4G_n, NET_290, VCC, SIM_RST);
    U74HC27 U10049(NET_300, NET_283, MDT11, R1C, GND, NET_303, GND, NET_301, NET_288, NET_287, NET_292, NET_297, NET_298, VCC, SIM_RST);
    U74LVC07 U10050(NET_229, __A10_2___CO_OUT, NET_301, __A10_2___RL1_n, NET_284, G11_n, GND, G11_n, NET_285, __A10_2___RL2_n, NET_216, __A10_2___L2_n, NET_255, VCC, SIM_RST);
    U74HC02 U10051(NET_289, L2GDG_n, __A10_1___L2_n, NET_286, WG1G_n, WL11_n, GND, G11_n, CGG, __A10_2___G1, RGG_n, G11_n, NET_292, VCC, SIM_RST);
    U74HC4002 U10052(NET_284, GND, SA11, NET_291, NET_290, NET_294, GND, NET_293, GND, SA12, NET_240, NET_239, NET_242, VCC, SIM_RST);
    wire U10053_3_NC;
    wire U10053_4_NC;
    wire U10053_5_NC;
    wire U10053_6_NC;
    wire U10053_8_NC;
    wire U10053_9_NC;
    wire U10053_10_NC;
    wire U10053_11_NC;
    U74HC27 #(1, 0, 0) U10053(NET_289, NET_286, U10053_3_NC, U10053_4_NC, U10053_5_NC, U10053_6_NC, GND, U10053_8_NC, U10053_9_NC, U10053_10_NC, U10053_11_NC, NET_285, __A10_2___G1, VCC, SIM_RST);
    U74HC02 U10054(NET_218, A2XG_n, __A10_2___A2_n, NET_232, WYLOG_n, WL12_n, GND, WL11_n, WYDG_n, NET_233, __A10_2__Y2_n, CUG, __A10_2__Y2, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U10055(MONEX, NET_218, __A10_2__X2_n, CLXC, CUG, __A10_2__X2, GND, __A10_2__Y2_n, NET_232, NET_233, __A10_2__Y2, __A10_2__X2_n, __A10_2__X2, VCC, SIM_RST);
    U74HC02 U10056(NET_230, __A10_2__X2_n, __A10_2__Y2_n, __A10_2___XUY2, __A10_2__X2, __A10_2__Y2, GND, XUY14_n, __A10_2___XUY2, NET_229, NET_230, __A10_2___XUY2, NET_228, VCC, SIM_RST);
    U74HC27 U10057(NET_230, __A10_2___XUY2, NET_230, __A10_2___SUMA2, __A10_2___CO_IN, __A10_2___CI_OUT, GND, NET_231, __A10_2___SUMA2, __A10_2___SUMB2, RULOG_n, __A10_2___SUMA2, __A10_2___CI_INTERNAL, VCC, SIM_RST);
    U74HC02 U10058(__A10_2___SUMB2, NET_228, NET_227, NET_217, WAG_n, WL12_n, GND, WL14_n, WALSG_n, NET_219, __A10_2___A2_n, CAG, NET_215, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U10059(NET_217, NET_219, NET_231, NET_214, CH12, NET_216, GND, NET_255, NET_258, NET_259, NET_251, __A10_2___A2_n, NET_215, VCC, SIM_RST);
    U74HC02 U10060(NET_214, RAG_n, __A10_2___A2_n, NET_258, WLG_n, WL12_n, GND, G15_n, G2LSG_n, NET_259, __A10_2___L2_n, CLG1G, NET_251, VCC, SIM_RST);
    U74HC27 U10061(RLG_n, __A10_2___L2_n, NET_253, NET_252, NET_220, NET_221, GND, NET_224, MDT12, R1C, GND, NET_253, GND, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U10062(NET_249, WQG_n, WL12_n, __A10_2___Q2_n, NET_249, NET_250, GND, __A10_2___Q2_n, CQG, NET_250, RQG_n, __A10_2___Q2_n, NET_252, VCC, SIM_RST);
    U74LVC07 U10063(NET_221, __A10_2___RL2_n, NET_222, __A10_2___Z2_n, NET_224, __A10_2___RL2_n, GND, __A10_2___RL2_n, NET_245, __A10_2___G2_n, NET_242, __A10_2___G2_n, NET_241, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U10064(NET_254, WZG_n, WL12_n, NET_222, NET_254, NET_223, GND, __A10_2___Z2_n, CZG, NET_223, RZG_n, __A10_2___Z2_n, NET_220, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U10065(NET_256, WBG_n, WL12_n, __A10_2___B2_n, NET_256, NET_257, GND, __A10_2___B2_n, CBG, NET_257, RBHG_n, __A10_2___B2_n, NET_244, VCC, SIM_RST);
    wire U10066_8_NC;
    wire U10066_9_NC;
    wire U10066_10_NC;
    wire U10066_11_NC;
    U74HC27 #(0, 1, 0) U10066(NET_244, NET_243, NET_238, NET_237, __A10_2___G2, NET_241, GND, U10066_8_NC, U10066_9_NC, U10066_10_NC, U10066_11_NC, NET_245, NET_248, VCC, SIM_RST);
    U74HC02 U10067(NET_243, NET_257, RCG_n, NET_240, WL11_n, WG3G_n, GND, WL13_n, WG4G_n, NET_239, L2GDG_n, __A10_2___L1_n, NET_238, VCC, SIM_RST);
    wire U10068_11_NC;
    wire U10068_12_NC;
    wire U10068_13_NC;
    U74HC02 U10068(NET_237, WG1G_n, WL12_n, __A10_2___G2, __A10_2___G2_n, CGG, GND, RGG_n, __A10_2___G2_n, NET_248, U10068_11_NC, U10068_12_NC, U10068_13_NC, VCC, SIM_RST);
    wire U10069_10_NC;
    wire U10069_11_NC;
    wire U10069_12_NC;
    wire U10069_13_NC;
    U74HC04 U10069(__A10_2___G2_n, __A10_2___GEM2, __A10_2___RL2_n, __A10_2___WL2, __A10_2___WL2, WL12_n, GND, __A10_2___MWL2, __A10_2___RL2_n, U10069_10_NC, U10069_11_NC, U10069_12_NC, U10069_13_NC, VCC, SIM_RST);
endmodule