`timescale 1ns/1ps
`default_nettype none

module counter_cell_ii(VCC, GND, SIM_RST, SIM_CLK, T12, T12A, INCSET_n, RSCT, BKTF_n, RSSB, BMAGXP, BMAGXM, BMAGYP, BMAGYM, EMSD, OTLNKM, ALTM, BMAGZP, BMAGZM, INLNKP, INLNKM, RNRADP, RNRADM, GYROD, XB0, XB1, XB2, XB3, XB4, XB5, XB6, XB7, OCTAD2, OCTAD3, OCTAD4, OCTAD5, OCTAD6, CG13, CG23, C24A, C25A, C26A, C27A, C30A, C31A, C32A, C32P, C32M, C33A, C33P, C33M, C34A, C34P, C34M, C35A, C35P, C35M, C36A, C36P, C36M, C37A, C37P, C37M, C40A, C40P, C40M, C41A, C41P, C41M, C50A, C51A, C52A, C53A, C54A, C55A, CA2_n, CA3_n, CA4_n, CA5_n, CA6_n, CXB0_n, CXB1_n, CXB2_n, CXB3_n, CXB4_n, CXB5_n, CXB6_n, CXB7_n, CAD1, CAD2, CAD3, CAD4, CAD5, CAD6, CG26, PINC, MINC, DINC, DINC_n, PCDU, MCDU, SHANC_n, SHIFT, SHIFT_n, CTROR, CTROR_n);
    input wire VCC;
    input wire GND;
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire ALTM;
    input wire BKTF_n;
    input wire BMAGXM;
    input wire BMAGXP;
    input wire BMAGYM;
    input wire BMAGYP;
    input wire BMAGZM;
    input wire BMAGZP;
    input wire C24A;
    input wire C25A;
    input wire C26A;
    input wire C27A;
    input wire C30A;
    input wire C31A;
    input wire C32A;
    input wire C32M;
    input wire C32P;
    input wire C33A;
    input wire C33M;
    input wire C33P;
    input wire C34A;
    input wire C34M;
    input wire C34P;
    input wire C35A;
    input wire C35M;
    input wire C35P;
    input wire C36A;
    input wire C36M;
    input wire C36P;
    input wire C37A;
    input wire C37M;
    input wire C37P;
    input wire C40A;
    input wire C40M;
    input wire C40P;
    input wire C41A;
    input wire C41M;
    input wire C41P;
    input wire C50A;
    input wire C51A;
    input wire C52A;
    input wire C53A;
    input wire C54A;
    input wire C55A;
    output wire CA2_n;
    output wire CA3_n;
    output wire CA4_n;
    output wire CA5_n;
    output wire CA6_n;
    output wire CAD1;
    output wire CAD2;
    output wire CAD3;
    output wire CAD4;
    output wire CAD5;
    output wire CAD6;
    input wire CG13;
    input wire CG23;
    output wire CG26;
    output wire CTROR;
    output wire CTROR_n;
    output wire CXB0_n;
    output wire CXB1_n;
    output wire CXB2_n;
    output wire CXB3_n;
    output wire CXB4_n;
    output wire CXB5_n;
    output wire CXB6_n;
    output wire CXB7_n;
    output wire DINC;
    output wire DINC_n;
    input wire EMSD;
    input wire GYROD;
    input wire INCSET_n;
    input wire INLNKM;
    input wire INLNKP;
    output wire MCDU;
    output wire MINC;
    input wire OCTAD2;
    input wire OCTAD3;
    input wire OCTAD4;
    input wire OCTAD5;
    input wire OCTAD6;
    input wire OTLNKM;
    output wire PCDU;
    output wire PINC;
    input wire RNRADM;
    input wire RNRADP;
    input wire RSCT;
    input wire RSSB;
    output wire SHANC_n;
    output wire SHIFT;
    output wire SHIFT_n;
    input wire T12;
    input wire T12A;
    input wire XB0;
    input wire XB1;
    input wire XB2;
    input wire XB3;
    input wire XB4;
    input wire XB5;
    input wire XB6;
    input wire XB7;
    wire __A21_1__30SUM;
    wire __A21_1__32004K; //FPGA#wand
    wire __A21_1__50SUM;
    wire __A21_1__C42A;
    wire __A21_1__C42M;
    wire __A21_1__C42P;
    wire __A21_1__C43A;
    wire __A21_1__C43M;
    wire __A21_1__C43P;
    wire __A21_1__C44A;
    wire __A21_1__C44M;
    wire __A21_1__C44P;
    wire __A21_1__C45A;
    wire __A21_1__C45M;
    wire __A21_1__C45P;
    wire __A21_1__C46A;
    wire __A21_1__C46M;
    wire __A21_1__C46P;
    wire __A21_1__C47A;
    wire __A21_1__C56A;
    wire __A21_1__C57A;
    wire __A21_1__C60A;
    wire __A21_1__DINCNC_n;
    wire __A21_1__MCDU_n;
    wire __A21_1__MINC_n;
    wire __A21_1__PCDU_n;
    wire __A21_1__PINC_n;
    wire __A21_1__RSCT_n;
    wire __A21_1__SHANC;
    wire __A21_1__SHINC;
    wire __A21_1__SHINC_n;
    wire __A21_3__C42R;
    wire __A21_3__C43R;
    wire __A21_3__C44R;
    wire __A21_3__C45R;
    wire __A21_3__C46R;
    wire __A21_3__C47R;
    wire __A21_3__C56R;
    wire __A21_3__C57R;
    wire __A21_3__C60R;
    wire __A21_3__CG15;
    wire __A21_3__CG16;
    wire __A21_NET_131;
    wire __A21_NET_132; //FPGA#wand
    wire __A21_NET_133;
    wire __A21_NET_137;
    wire __A21_NET_139;
    wire __A21_NET_140;
    wire __A21_NET_141; //FPGA#wand
    wire __A21_NET_142;
    wire __A21_NET_143;
    wire __A21_NET_144; //FPGA#wand
    wire __A21_NET_145; //FPGA#wand
    wire __A21_NET_146; //FPGA#wand
    wire __A21_NET_147;
    wire __A21_NET_148; //FPGA#wand
    wire __A21_NET_149;
    wire __A21_NET_151;
    wire __A21_NET_152;
    wire __A21_NET_153;
    wire __A21_NET_154;
    wire __A21_NET_156; //FPGA#wand
    wire __A21_NET_157;
    wire __A21_NET_158; //FPGA#wand
    wire __A21_NET_159;
    wire __A21_NET_160;
    wire __A21_NET_161;
    wire __A21_NET_162;
    wire __A21_NET_163;
    wire __A21_NET_166;
    wire __A21_NET_167;
    wire __A21_NET_168;
    wire __A21_NET_171;
    wire __A21_NET_172;
    wire __A21_NET_181;
    wire __A21_NET_182;
    wire __A21_NET_183;
    wire __A21_NET_188;
    wire __A21_NET_192;
    wire __A21_NET_197;
    wire __A21_NET_202;
    wire __A21_NET_203;
    wire __A21_NET_204; //FPGA#wand
    wire __A21_NET_205;
    wire __A21_NET_206;
    wire __A21_NET_208;
    wire __A21_NET_210;
    wire __A21_NET_211;
    wire __A21_NET_216;
    wire __A21_NET_219;
    wire __A21_NET_220;
    wire __A21_NET_221;
    wire __A21_NET_222; //FPGA#wand
    wire __A21_NET_227;
    wire __A21_NET_228; //FPGA#wand
    wire __A21_NET_229;
    wire __A21_NET_230;
    wire __A21_NET_231;
    wire __A21_NET_232;
    wire __A21_NET_233;
    wire __A21_NET_235;
    wire __A21_NET_236;
    wire __A21_NET_237;
    wire __A21_NET_238;
    wire __A21_NET_239;
    wire __A21_NET_240;
    wire __A21_NET_243;
    wire __A21_NET_244;
    wire __A21_NET_245;
    wire __A21_NET_246;
    wire __A21_NET_247;
    wire __A21_NET_248;
    wire __A21_NET_249;
    wire __A21_NET_251;
    wire __A21_NET_252;
    wire __A21_NET_253;
    wire __A21_NET_254;
    wire __A21_NET_256;
    wire __A21_NET_257;
    wire __A21_NET_258;
    wire __A21_NET_259;
    wire __A21_NET_260;
    wire __A21_NET_261;
    wire __A21_NET_263;
    wire __A21_NET_264;
    wire __A21_NET_265;
    wire __A21_NET_266;
    wire __A21_NET_267;
    wire __A21_NET_268;
    wire __A21_NET_269;
    wire __A21_NET_270;
    wire __A21_NET_271;
    wire __A21_NET_272;
    wire __A21_NET_273;
    wire __A21_NET_274;
    wire __A21_NET_275;
    wire __A21_NET_277;
    wire __A21_NET_278;
    wire __A21_NET_279;
    wire __A21_NET_280;
    wire __A21_NET_281;
    wire __A21_NET_282;
    wire __A21_NET_284;
    wire __A21_NET_285;
    wire __A21_NET_286;
    wire __A21_NET_287;
    wire __A21_NET_289;
    wire __A21_NET_290;
    wire __A21_NET_291;
    wire __A21_NET_294;
    wire __A21_NET_297;
    wire __A21_NET_298;
    wire __A21_NET_299;
    wire __A21_NET_300;
    wire __A21_NET_301;
    wire __A21_NET_302;
    wire __A21_NET_303;
    wire __A21_NET_304;
    wire __A21_NET_305;
    wire __A21_NET_306;
    wire __A21_NET_309;
    wire __A21_NET_310;
    wire __A21_NET_311;

    pullup R21001(__A21_NET_204);
    pullup R21002(__A21_NET_146);
    pullup R21003(__A21_NET_145);
    pullup R21004(__A21_1__32004K);
    pullup R21005(__A21_NET_148);
    pullup R21006(__A21_NET_144);
    pullup R21007(__A21_NET_222);
    pullup R21008(__A21_NET_228);
    pullup R21009(__A21_NET_132);
    pullup R21010(__A21_NET_141);
    pullup R21011(__A21_NET_156);
    pullup R21012(__A21_NET_158);
    U74HC4002 U21001(__A21_NET_203, C25A, C27A, C31A, C33A,  , GND,  , C35A, C37A, C41A, __A21_1__C43A, __A21_NET_202, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U21002(__A21_NET_203, __A21_NET_204, __A21_NET_202, __A21_NET_204, __A21_NET_192, __A21_NET_204, GND, __A21_NET_204, __A21_NET_197, __A21_NET_146, __A21_NET_211, __A21_NET_146, __A21_NET_210, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC4002 U21003(__A21_NET_192, __A21_1__C45A, __A21_1__C47A, C51A, C53A,  , GND,  , C26A, C27A, C32A, C33A, __A21_NET_211, VCC, SIM_RST, SIM_CLK);
    U74HC02 U21004(__A21_NET_197, C55A, __A21_1__C57A, __A21_NET_205, __A21_1__C56A, __A21_1__C57A, GND, __A21_1__30SUM, __A21_1__C60A, __A21_NET_221, __A21_1__50SUM, __A21_1__C60A, __A21_NET_219, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21005(__A21_NET_210, C36A, C37A, __A21_1__C42A, __A21_1__C43A,  , GND,  , __A21_1__C46A, __A21_1__C47A, C52A, C53A, __A21_NET_206, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U21006(__A21_NET_206, __A21_NET_146, __A21_NET_205, __A21_NET_146, __A21_NET_208, __A21_NET_145, GND, __A21_NET_145, __A21_NET_171, __A21_NET_145, __A21_NET_172, __A21_NET_145, __A21_NET_167, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC4002 U21007(__A21_NET_208, C24A, C25A, C26A, C27A,  , GND,  , C34A, C35A, C36A, C37A, __A21_NET_171, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21008(__A21_NET_172, __A21_1__C44A, __A21_1__C45A, __A21_1__C46A, __A21_1__C47A,  , GND,  , C54A, C55A, __A21_1__C56A, __A21_1__C57A, __A21_NET_167, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21009(__A21_NET_166, C30A, C31A, C32A, C33A,  , GND,  , C34A, C35A, C36A, C37A, __A21_NET_168, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U21010(__A21_NET_166, __A21_1__32004K, __A21_NET_168, __A21_1__32004K, __A21_NET_188, __A21_NET_148, GND, __A21_NET_148, __A21_NET_182, __A21_NET_144, __A21_NET_181, __A21_NET_144, __A21_NET_221, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC04 U21011(__A21_1__32004K, __A21_1__30SUM, __A21_NET_148, __A21_1__50SUM, DINC, DINC_n, GND, CXB0_n, XB0, CXB1_n, XB1, CXB2_n, XB2, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21012(__A21_NET_188, C50A, C51A, C52A, C53A,  , GND,  , C54A, C55A, __A21_1__C56A, __A21_1__C57A, __A21_NET_182, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21013(__A21_NET_181, C24A, C25A, C26A, C27A,  , GND,  , C40A, C41A, __A21_1__C42A, __A21_1__C43A, __A21_NET_183, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U21015(__A21_NET_183, __A21_NET_222, __A21_NET_220, __A21_NET_222, __A21_NET_219, __A21_NET_222, GND, __A21_NET_228, __A21_NET_229, __A21_NET_228, __A21_NET_227, __A21_NET_228, __A21_NET_216, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC4002 U21016(__A21_NET_220, __A21_1__C44A, __A21_1__C45A, __A21_1__C46A, __A21_1__C47A,  , GND,  , __A21_1__C45M, __A21_1__C46M, __A21_1__C57A, __A21_1__C60A, __A21_NET_152, VCC, SIM_RST, SIM_CLK);
    U74HC02 U21017(__A21_NET_147, __A21_1__30SUM, __A21_1__50SUM, CAD1, __A21_1__RSCT_n, __A21_NET_204, GND, __A21_1__RSCT_n, __A21_NET_146, CAD2, __A21_1__RSCT_n, __A21_NET_145, CAD3, VCC, SIM_RST, SIM_CLK);
    U74HC02 U21018(CAD4, __A21_1__RSCT_n, __A21_NET_147, CAD5, __A21_1__RSCT_n, __A21_NET_144, GND, __A21_1__RSCT_n, __A21_NET_222, CAD6, __A21_1__C45P, __A21_1__C46P, __A21_NET_151, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21019(C31A, __A21_1__C47A, C51A, C52A, C53A, __A21_NET_227, GND, __A21_NET_216, C54A, C55A, __A21_1__C56A, __A21_NET_229, C50A, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U21020(__A21_NET_154, INCSET_n, __A21_NET_152, __A21_NET_153, INCSET_n, __A21_NET_151, GND, INCSET_n, __A21_NET_228, __A21_NET_149, __A21_NET_154, __A21_1__SHINC, __A21_1__SHINC_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21021(__A21_1__SHINC, __A21_1__SHINC_n, T12A, SHANC_n, __A21_NET_153, __A21_1__SHANC, GND, SHANC_n, T12A, __A21_1__SHANC, __A21_NET_149, DINC, __A21_1__DINCNC_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U21022(DINC, __A21_1__DINCNC_n, T12A, __A21_NET_131, INCSET_n, __A21_NET_132, GND, __A21_NET_131, PINC, __A21_1__PINC_n, __A21_1__PINC_n, T12, PINC, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21023(__A21_NET_133, C24A, C25A, C26A, C27A,  , GND,  , C30A, C37P, C40P, C41P, __A21_NET_137, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U21024(__A21_NET_133, __A21_NET_132, __A21_NET_137, __A21_NET_132, __A21_NET_143, __A21_NET_132, GND, __A21_NET_141, __A21_NET_140, __A21_NET_141, __A21_NET_139, __A21_NET_156, __A21_NET_160, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 U21025(__A21_1__C42P, __A21_1__C43P, __A21_1__C42M, __A21_1__C43M, __A21_1__C44M, __A21_NET_140, GND, __A21_NET_139, C37M, C40M, C41M, __A21_NET_143, __A21_1__C44P, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21026(__A21_NET_142, INCSET_n, __A21_NET_141, __A21_1__MINC_n, __A21_NET_142, MINC, GND, __A21_1__MINC_n, T12A, MINC, C35P, C36P, __A21_NET_157, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21027(C32P, C33P, C32M, C33M, C34M, __A21_NET_159, GND,  ,  ,  ,  , __A21_NET_160, C34P, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U21028(__A21_NET_157, __A21_NET_156, __A21_NET_159, __A21_NET_158, __A21_NET_163, __A21_NET_158, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21029(__A21_NET_161, INCSET_n, __A21_NET_156, __A21_1__PCDU_n, __A21_NET_161, PCDU, GND, __A21_1__PCDU_n, T12A, PCDU, C35M, C36M, __A21_NET_163, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21030(__A21_NET_162, INCSET_n, __A21_NET_158, __A21_1__MCDU_n, __A21_NET_162, MCDU, GND, __A21_1__MCDU_n, T12A, MCDU,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21031(__A21_NET_284, BMAGXP, __A21_NET_282, __A21_NET_282, __A21_NET_284, __A21_3__C42R, GND, BMAGXM, __A21_NET_279, __A21_NET_285, __A21_NET_285, __A21_3__C42R, __A21_NET_279, VCC, SIM_RST, SIM_CLK);
    U74HC04 U21032(BKTF_n, __A21_NET_270, RSSB, __A21_NET_306, __A21_NET_303, __A21_3__CG15, GND, CTROR, CTROR_n, __A21_NET_240, RSSB, __A21_NET_238, BKTF_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21033(__A21_NET_280, __A21_NET_282, __A21_NET_279, __A21_NET_281, __A21_NET_270, __A21_NET_280, GND, __A21_NET_281, __A21_NET_302, __A21_NET_286, __A21_NET_286, __A21_3__C42R, __A21_NET_302, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21034(__A21_1__C42A, CG13, __A21_NET_286, __A21_NET_275, BMAGYP, __A21_NET_273, GND, __A21_1__SHINC, __A21_1__SHANC, SHIFT_n, BMAGYM, __A21_NET_272, __A21_NET_274, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21035(__A21_NET_306, CA4_n, __A21_NET_284, CA4_n, CXB2_n, __A21_1__C42P, GND, __A21_1__C42M, __A21_NET_285, CA4_n, CXB2_n, __A21_3__C42R, CXB2_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21036(__A21_NET_272, __A21_NET_274, __A21_3__C43R, __A21_NET_269, __A21_NET_273, __A21_NET_272, GND, __A21_NET_270, __A21_NET_269, __A21_NET_271, __A21_NET_271, __A21_NET_278, __A21_NET_277, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21037(__A21_NET_278, __A21_NET_277, __A21_3__C43R, __A21_NET_300, EMSD, __A21_NET_301, GND, __A21_NET_300, __A21_3__C56R, __A21_NET_301, __A21_NET_270, __A21_NET_300, __A21_NET_311, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21038(__A21_NET_306, CA4_n, __A21_NET_275, CA4_n, CXB3_n, __A21_1__C43P, GND, __A21_1__C43M, __A21_NET_274, CA4_n, CXB3_n, __A21_3__C43R, CXB3_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21039(CG13, __A21_NET_302, CG13, __A21_NET_302, __A21_NET_278, __A21_NET_303, GND, __A21_3__C56R, __A21_NET_306, CA5_n, CXB6_n, __A21_1__C43A, __A21_NET_277, VCC, SIM_RST, SIM_CLK);
    U74HC02 U2104( ,  ,  ,  ,  ,  , GND, __A21_NET_275, __A21_3__C43R, __A21_NET_273,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U21040(__A21_NET_309, __A21_NET_311, __A21_NET_310, __A21_NET_310, __A21_NET_309, __A21_3__C56R, GND, CG23, __A21_NET_309, __A21_1__C56A, OTLNKM, __A21_NET_304, __A21_NET_305, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U21041(__A21_NET_304, __A21_NET_305, __A21_3__C57R, __A21_NET_290, __A21_NET_270, __A21_NET_305, GND, __A21_NET_290, __A21_NET_294, __A21_NET_291, __A21_NET_291, __A21_3__C57R, __A21_NET_294, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21042(__A21_NET_306, CA5_n, CG23, __A21_NET_310, __A21_NET_291, __A21_1__C57A, GND, __A21_3__C60R, __A21_NET_306, CA6_n, CXB0_n, __A21_3__C57R, CXB7_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U21043(__A21_NET_289, ALTM, __A21_NET_287, __A21_NET_287, __A21_NET_289, __A21_3__C60R, GND, __A21_NET_270, __A21_NET_289, __A21_NET_297, __A21_NET_297, __A21_NET_299, __A21_NET_298, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21044(__A21_NET_299, __A21_NET_298, __A21_3__C60R, __A21_NET_247, BMAGZP, __A21_NET_246, GND, __A21_NET_247, __A21_3__C44R, __A21_NET_246, BMAGZM, __A21_NET_244, __A21_NET_243, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21045(__A21_1__C60A, CG23, __A21_NET_310, __A21_NET_294, __A21_NET_298,  , GND,  , CG23, __A21_NET_310, __A21_NET_294, __A21_NET_299, CTROR_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21046(__A21_NET_244, __A21_NET_243, __A21_3__C44R, __A21_NET_245, __A21_NET_246, __A21_NET_244, GND, __A21_NET_238, __A21_NET_245, __A21_NET_249, __A21_NET_249, __A21_NET_263, __A21_NET_248, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U21047(__A21_NET_263, __A21_NET_248, __A21_3__C44R, __A21_1__C44A, __A21_3__CG15, __A21_NET_248, GND, INLNKP, __A21_NET_232, __A21_NET_233, __A21_NET_233, __A21_3__C45R, __A21_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21048(__A21_NET_240, CA4_n, __A21_NET_247, CA4_n, CXB4_n, __A21_1__C44P, GND, __A21_1__C44M, __A21_NET_243, CA4_n, CXB4_n, __A21_3__C44R, CXB4_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21049(__A21_NET_235, INLNKM, __A21_NET_230, __A21_NET_230, __A21_NET_235, __A21_3__C45R, GND, __A21_NET_232, __A21_NET_230, __A21_NET_231, __A21_NET_238, __A21_NET_231, __A21_NET_239, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21050(__A21_NET_237, __A21_NET_239, __A21_NET_236, __A21_NET_236, __A21_NET_237, __A21_3__C45R, GND, RNRADP, __A21_NET_260, __A21_NET_259, __A21_NET_259, __A21_3__C46R, __A21_NET_260, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21051(__A21_NET_240, CA4_n, __A21_NET_233, CA4_n, CXB5_n, __A21_1__C45P, GND, __A21_1__C45M, __A21_NET_235, CA4_n, CXB5_n, __A21_3__C45R, CXB5_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21052(__A21_3__CG15, __A21_NET_263, __A21_3__CG15, __A21_NET_263, __A21_NET_236, __A21_NET_261, GND, __A21_3__C46R, __A21_NET_240, CA4_n, CXB6_n, __A21_1__C45A, __A21_NET_237, VCC, SIM_RST, SIM_CLK);
    U74HC04 U21053(__A21_NET_261, __A21_3__CG16, __A21_NET_257, CG26, XB3, CXB3_n, GND, CXB4_n, XB4, CXB5_n, XB5, CXB6_n, XB6, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21054(__A21_NET_267, __A21_NET_238, __A21_NET_258, __A21_NET_268, __A21_NET_267, __A21_NET_266, GND, __A21_NET_268, __A21_3__C46R, __A21_NET_266, __A21_3__CG16, __A21_NET_268, __A21_1__C46A, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21055(__A21_NET_265, RNRADM, __A21_NET_264, __A21_NET_264, __A21_NET_265, __A21_3__C46R, GND, __A21_NET_260, __A21_NET_264, __A21_NET_258,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21056( ,  ,  , __A21_NET_253, GYROD, __A21_NET_254, GND, __A21_NET_253, __A21_3__C47R, __A21_NET_254, __A21_NET_238, __A21_NET_253, __A21_NET_252, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21057(__A21_NET_259, CA4_n, CA4_n, CXB6_n, __A21_NET_265, __A21_1__C46M, GND, __A21_3__C47R, __A21_NET_240, CA4_n, CXB7_n, __A21_1__C46P, CXB6_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U21058(__A21_NET_251, __A21_NET_252, __A21_NET_256, __A21_NET_256, __A21_NET_251, __A21_3__C47R, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U21059(__A21_3__CG16, __A21_NET_266, __A21_3__CG16, __A21_NET_266, __A21_NET_256, __A21_NET_257, GND,  ,  ,  ,  , __A21_1__C47A, __A21_NET_251, VCC, SIM_RST, SIM_CLK);
    U74HC04 U21060(XB7, CXB7_n, OCTAD2, CA2_n, OCTAD3, CA3_n, GND, CA4_n, OCTAD4, CA5_n, OCTAD5, CA6_n, OCTAD6, VCC, SIM_RST, SIM_CLK);
    U74HC04 U21061(SHIFT_n, SHIFT, RSCT, __A21_1__RSCT_n,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
endmodule