`timescale 1ns/1ps

module four_bit_1(VCC, GND, SIM_RST, A2XG_n, CAG, CBG, CGG, CLG1G, CLXC, CQG, CUG, CZG, L2GDG_n, RAG_n, RCG_n, RGG_n, RLG_n, RQG_n, RZG_n, WAG_n, WALSG_n, WBG_n, WLG_n, WQG_n, WZG_n, CI01_n, MONEX, PONEX, TWOX, XUY05_n, XUY06_n, CH01, CH02, CH03, CH04, G01ED, G02ED, G03ED, G04ED, MCRO_n, G2LSG_n, G05_n, G06_n, G07_n, MDT01, MDT02, MDT03, MDT04, SA01, SA02, SA03, SA04, RBLG_n, RULOG_n, WL05_n, WL06_n, WG1G_n, WG3G_n, WG4G_n, WYDLOG_n, WYDG_n, WYLOG_n, RB1, R1C, R15, RB2, WL16_n, WHOMP, WHOMPA, CI05_n, CO06, G01, G01_n, G02, G03, G04, L01_n, L02_n, L04_n, WL01_n, WL02_n, WL03_n, WL04_n, XUY01_n, XUY02_n);
    input wire SIM_RST;
    input wire A2XG_n;
    input wire CAG;
    input wire CBG;
    input wire CGG;
    input wire CH01;
    input wire CH02;
    input wire CH03;
    input wire CH04;
    input wire CI01_n;
    output wire CI05_n;
    input wire CLG1G;
    input wire CLXC;
    inout wire CO06;
    input wire CQG;
    input wire CUG;
    input wire CZG;
    output wire G01;
    input wire G01ED;
    inout wire G01_n;
    output wire G02;
    input wire G02ED;
    output wire G03;
    input wire G03ED;
    output wire G04;
    input wire G04ED;
    input wire G05_n;
    input wire G06_n;
    input wire G07_n;
    input wire G2LSG_n;
    input wire GND;
    inout wire L01_n;
    inout wire L02_n;
    inout wire L04_n;
    input wire L2GDG_n;
    input wire MCRO_n;
    input wire MDT01;
    input wire MDT02;
    input wire MDT03;
    input wire MDT04;
    input wire MONEX;
    wire NET_137;
    wire NET_138;
    wire NET_139;
    wire NET_140;
    wire NET_141;
    wire NET_142;
    wire NET_143;
    wire NET_144;
    wire NET_145;
    wire NET_146;
    wire NET_147;
    wire NET_148;
    wire NET_149;
    wire NET_152;
    wire NET_155;
    wire NET_156;
    wire NET_157;
    wire NET_158;
    wire NET_159;
    wire NET_160;
    wire NET_161;
    wire NET_162;
    wire NET_163;
    wire NET_164;
    wire NET_167;
    wire NET_168;
    wire NET_169;
    wire NET_170;
    wire NET_173;
    wire NET_174;
    wire NET_175;
    wire NET_176;
    wire NET_177;
    wire NET_178;
    wire NET_179;
    wire NET_180;
    wire NET_181;
    wire NET_182;
    wire NET_183;
    wire NET_184;
    wire NET_185;
    wire NET_186;
    wire NET_187;
    wire NET_188;
    wire NET_189;
    wire NET_190;
    wire NET_191;
    wire NET_192;
    wire NET_193;
    wire NET_194;
    wire NET_195;
    wire NET_196;
    wire NET_197;
    wire NET_198;
    wire NET_199;
    wire NET_200;
    wire NET_205;
    wire NET_206;
    wire NET_207;
    wire NET_209;
    wire NET_210;
    wire NET_211;
    wire NET_212;
    wire NET_213;
    wire NET_214;
    wire NET_215;
    wire NET_216;
    wire NET_217;
    wire NET_218;
    wire NET_219;
    wire NET_220;
    wire NET_221;
    wire NET_222;
    wire NET_223;
    wire NET_224;
    wire NET_225;
    wire NET_226;
    wire NET_227;
    wire NET_228;
    wire NET_229;
    wire NET_230;
    wire NET_231;
    wire NET_232;
    wire NET_233;
    wire NET_234;
    wire NET_235;
    wire NET_236;
    wire NET_237;
    wire NET_238;
    wire NET_239;
    wire NET_240;
    wire NET_241;
    wire NET_242;
    wire NET_245;
    wire NET_248;
    wire NET_249;
    wire NET_250;
    wire NET_251;
    wire NET_252;
    wire NET_253;
    wire NET_254;
    wire NET_255;
    wire NET_256;
    wire NET_257;
    wire NET_260;
    wire NET_261;
    wire NET_262;
    wire NET_263;
    wire NET_266;
    wire NET_267;
    wire NET_268;
    wire NET_269;
    wire NET_270;
    wire NET_271;
    wire NET_272;
    wire NET_273;
    wire NET_274;
    wire NET_275;
    wire NET_276;
    wire NET_277;
    wire NET_278;
    wire NET_279;
    wire NET_280;
    wire NET_281;
    wire NET_282;
    wire NET_283;
    wire NET_284;
    wire NET_285;
    wire NET_286;
    wire NET_287;
    wire NET_288;
    wire NET_289;
    wire NET_290;
    wire NET_291;
    wire NET_293;
    wire NET_294;
    wire NET_298;
    wire NET_299;
    wire NET_300;
    wire NET_302;
    wire NET_303;
    wire NET_304;
    wire NET_305;
    wire NET_306;
    wire NET_307;
    wire NET_308;
    wire NET_309;
    wire NET_310;
    wire NET_311;
    wire NET_312;
    wire NET_313;
    wire NET_314;
    wire NET_315;
    wire NET_316;
    wire NET_317;
    wire NET_318;
    wire NET_319;
    wire NET_320;
    wire NET_321;
    wire NET_322;
    input wire PONEX;
    input wire R15;
    input wire R1C;
    input wire RAG_n;
    input wire RB1;
    input wire RB2;
    input wire RBLG_n;
    input wire RCG_n;
    input wire RGG_n;
    input wire RLG_n;
    input wire RQG_n;
    input wire RULOG_n;
    input wire RZG_n;
    input wire SA01;
    input wire SA02;
    input wire SA03;
    input wire SA04;
    input wire TWOX;
    input wire VCC;
    input wire WAG_n;
    input wire WALSG_n;
    input wire WBG_n;
    input wire WG1G_n;
    input wire WG3G_n;
    input wire WG4G_n;
    input wire WHOMP;
    input wire WHOMPA;
    output wire WL01_n;
    output wire WL02_n;
    output wire WL03_n;
    output wire WL04_n;
    input wire WL05_n;
    input wire WL06_n;
    input wire WL16_n;
    input wire WLG_n;
    input wire WQG_n;
    input wire WYDG_n;
    input wire WYDLOG_n;
    input wire WYLOG_n;
    input wire WZG_n;
    output wire XUY01_n;
    output wire XUY02_n;
    input wire XUY05_n;
    input wire XUY06_n;
    wire __A08_1__X1;
    wire __A08_1__X1_n;
    wire __A08_1__X2;
    wire __A08_1__X2_n;
    wire __A08_1__Y1;
    wire __A08_1__Y1_n;
    wire __A08_1__Y2;
    wire __A08_1__Y2_n;
    wire __A08_1___A1_n;
    wire __A08_1___A2_n;
    wire __A08_1___B1_n;
    wire __A08_1___B2_n;
    wire __A08_1___CI_INTERNAL;
    wire __A08_1___G2_n;
    wire __A08_1___GEM1;
    wire __A08_1___GEM2;
    wire __A08_1___MWL1;
    wire __A08_1___MWL2;
    wire __A08_1___Q1_n;
    wire __A08_1___Q2_n;
    wire __A08_1___RL1_n;
    wire __A08_1___RL2_n;
    wire __A08_1___RL_OUT_1;
    wire __A08_1___RL_OUT_2;
    wire __A08_1___SUMA1;
    wire __A08_1___SUMA2;
    wire __A08_1___SUMB1;
    wire __A08_1___SUMB2;
    wire __A08_1___WL1;
    wire __A08_1___WL2;
    wire __A08_1___Z1_n;
    wire __A08_1___Z2_n;
    wire __A08_2__X1;
    wire __A08_2__X1_n;
    wire __A08_2__X2;
    wire __A08_2__X2_n;
    wire __A08_2__Y1;
    wire __A08_2__Y1_n;
    wire __A08_2__Y2;
    wire __A08_2__Y2_n;
    wire __A08_2___A1_n;
    wire __A08_2___A2_n;
    wire __A08_2___B1_n;
    wire __A08_2___B2_n;
    wire __A08_2___CI_IN;
    wire __A08_2___CI_INTERNAL;
    wire __A08_2___CO_IN;
    wire __A08_2___G1_n;
    wire __A08_2___G2_n;
    wire __A08_2___GEM1;
    wire __A08_2___GEM2;
    wire __A08_2___L1_n;
    wire __A08_2___MWL1;
    wire __A08_2___MWL2;
    wire __A08_2___Q1_n;
    wire __A08_2___Q2_n;
    wire __A08_2___RL1_n;
    wire __A08_2___RL2_n;
    wire __A08_2___RL_OUT_1;
    wire __A08_2___RL_OUT_2;
    wire __A08_2___SUMA1;
    wire __A08_2___SUMA2;
    wire __A08_2___SUMB1;
    wire __A08_2___SUMB2;
    wire __A08_2___WL1;
    wire __A08_2___WL2;
    wire __A08_2___XUY1;
    wire __A08_2___XUY2;
    wire __A08_2___Z1_n;
    wire __A08_2___Z2_n;

    pullup R8001(__A08_2___CO_IN);
    pullup R8002(__A08_1___RL1_n);
    pullup R8003(L01_n);
    pullup R8005(__A08_1___Z1_n);
    pullup R8006(G01_n);
    pullup R8007(__A08_1___RL2_n);
    pullup R8008(L02_n);
    pullup R8009(__A08_1___Z2_n);
    pullup R8010(__A08_1___G2_n);
    pullup R8011(CO06);
    pullup R8012(__A08_2___RL1_n);
    pullup R8013(__A08_2___L1_n);
    pullup R8015(__A08_2___Z1_n);
    pullup R8016(__A08_2___G1_n);
    pullup R8017(__A08_2___RL2_n);
    pullup R8018(L04_n);
    pullup R8019(__A08_2___Z2_n);
    pullup R8020(__A08_2___G2_n);
    U74HC02 U8001(NET_205, A2XG_n, __A08_1___A1_n, NET_200, WYLOG_n, WL01_n, GND, WL16_n, WYDLOG_n, NET_199, __A08_1__Y1_n, CUG, __A08_1__Y1, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U8002(PONEX, NET_205, __A08_1__X1_n, CLXC, CUG, __A08_1__X1, GND, __A08_1__Y1_n, NET_200, NET_199, __A08_1__Y1, __A08_1__X1_n, __A08_1__X1, VCC, SIM_RST);
    U74HC02 U8003(NET_209, __A08_1__X1_n, __A08_1__Y1_n, XUY01_n, __A08_1__X1, __A08_1__Y1, GND, NET_209, XUY01_n, NET_207, NET_209, __A08_1___SUMA1, __A08_1___CI_INTERNAL, VCC, SIM_RST);
    wire U8004_1_NC;
    wire U8004_2_NC;
    wire U8004_12_NC;
    wire U8004_13_NC;
    U74HC27 U8004(U8004_1_NC, U8004_2_NC, __A08_1___SUMA1, __A08_1___SUMB1, RULOG_n, NET_187, GND, NET_191, __A08_2___XUY1, XUY01_n, CI01_n, U8004_12_NC, U8004_13_NC, VCC, SIM_RST);
    U74HC04 U8005(CI01_n, NET_206, G01_n, __A08_1___GEM1, __A08_1___RL1_n, __A08_1___WL1, GND, WL01_n, __A08_1___WL1, __A08_1___MWL1, __A08_1___RL1_n, NET_157, __A08_1___CI_INTERNAL, VCC, SIM_RST);
    U74HC02 U8006(__A08_1___SUMB1, NET_207, NET_206, NET_190, WAG_n, WL01_n, GND, WL03_n, WALSG_n, NET_192, __A08_1___A1_n, CAG, NET_188, VCC, SIM_RST);
    U74LVC07 U8007(NET_191, __A08_2___CO_IN, NET_185, __A08_1___RL1_n, NET_198, L01_n, GND, __A08_1___Z1_n, NET_221, __A08_1___RL1_n, NET_222, __A08_1___RL1_n, NET_220, VCC, SIM_RST);
    U74HC02 U8008(NET_186, RAG_n, __A08_1___A1_n, NET_189, WLG_n, WL01_n, GND, __A08_2___G2_n, G2LSG_n, NET_196, L01_n, CLG1G, NET_197, VCC, SIM_RST);
    wire U8009_1_NC;
    wire U8009_2_NC;
    wire U8009_3_NC;
    U74HC02 #(0, 0, 1, 0) U8009(U8009_1_NC, U8009_2_NC, U8009_3_NC, NET_194, WQG_n, WL01_n, GND, NET_194, NET_193, __A08_1___Q1_n, __A08_1___Q1_n, CQG, NET_193, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U8010(NET_195, RQG_n, __A08_1___Q1_n, NET_224, WZG_n, WL01_n, GND, NET_224, NET_223, NET_221, __A08_1___Z1_n, CZG, NET_223, VCC, SIM_RST);
    U74HC27 U8011(__A08_1___RL_OUT_1, NET_195, MDT01, RB1, R15, NET_220, GND, NET_227, NET_225, NET_226, NET_212, NET_222, NET_219, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U8012(NET_219, RZG_n, __A08_1___Z1_n, NET_228, WBG_n, WL01_n, GND, NET_228, NET_229, __A08_1___B1_n, __A08_1___B1_n, CBG, NET_229, VCC, SIM_RST);
    U74LVC07 U8013(NET_170, __A08_2___CO_IN, NET_227, __A08_1___RL1_n, NET_211, G01_n, GND, G01_n, NET_210, __A08_1___RL2_n, NET_137, L02_n, NET_147, VCC, SIM_RST);
    U74HC02 U8014(NET_225, RBLG_n, __A08_1___B1_n, NET_226, NET_229, RCG_n, GND, WL16_n, WG3G_n, NET_216, WL02_n, WG4G_n, NET_215, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U8015(NET_190, NET_192, NET_187, NET_186, CH01, NET_185, GND, NET_198, NET_189, NET_196, NET_197, __A08_1___A1_n, NET_188, VCC, SIM_RST);
    U74HC02 U8016(NET_214, L2GDG_n, MCRO_n, NET_213, WG1G_n, WL01_n, GND, G01_n, CGG, G01, RGG_n, G01_n, NET_212, VCC, SIM_RST);
    U74HC27 #(1, 0, 0) U8017(NET_214, NET_213, WHOMPA, __A08_2___XUY2, XUY02_n, NET_170, GND, __A08_1___RL_OUT_1, RLG_n, L01_n, GND, NET_210, G01, VCC, SIM_RST);
    U74HC4002 #(1, 0) U8018(NET_211, G01ED, SA01, NET_216, NET_215, NET_218, GND, NET_217, G02ED, SA02, NET_164, NET_163, NET_162, VCC, SIM_RST);
    U74HC02 U8019(NET_158, A2XG_n, __A08_1___A2_n, NET_160, WYLOG_n, WL02_n, GND, WL01_n, WYDG_n, NET_159, __A08_1__Y2_n, CUG, __A08_1__Y2, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U8020(TWOX, NET_158, __A08_1__X2_n, CLXC, CUG, __A08_1__X2, GND, __A08_1__Y2_n, NET_160, NET_159, __A08_1__Y2, __A08_1__X2_n, __A08_1__X2, VCC, SIM_RST);
    wire U8021_8_NC;
    wire U8021_9_NC;
    wire U8021_10_NC;
    U74HC02 U8021(NET_152, __A08_1__X2_n, __A08_1__Y2_n, XUY02_n, __A08_1__X2, __A08_1__Y2, GND, U8021_8_NC, U8021_9_NC, U8021_10_NC, NET_152, XUY02_n, NET_155, VCC, SIM_RST);
    wire U8022_1_NC;
    wire U8022_2_NC;
    wire U8022_12_NC;
    wire U8022_13_NC;
    U74HC27 U8022(U8022_1_NC, U8022_2_NC, NET_152, __A08_1___SUMA2, GND, __A08_2___CI_IN, GND, NET_156, __A08_1___SUMA2, __A08_1___SUMB2, RULOG_n, U8022_12_NC, U8022_13_NC, VCC, SIM_RST);
    U74HC02 U8023(__A08_1___SUMB2, NET_155, NET_157, NET_141, WAG_n, WL02_n, GND, WL04_n, WALSG_n, NET_140, __A08_1___A2_n, CAG, NET_139, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U8024(NET_141, NET_140, NET_156, NET_142, CH02, NET_137, GND, NET_147, NET_175, NET_176, NET_177, __A08_1___A2_n, NET_139, VCC, SIM_RST);
    U74HC02 U8025(NET_142, RAG_n, __A08_1___A2_n, NET_175, WLG_n, WL02_n, GND, G05_n, G2LSG_n, NET_176, L02_n, CLG1G, NET_177, VCC, SIM_RST);
    U74HC27 U8026(RLG_n, L02_n, __A08_1___RL_OUT_2, NET_143, NET_149, NET_148, GND, NET_138, MDT02, R1C, RB2, __A08_1___RL_OUT_2, GND, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U8027(NET_179, WQG_n, WL02_n, __A08_1___Q2_n, NET_179, NET_178, GND, __A08_1___Q2_n, CQG, NET_178, RQG_n, __A08_1___Q2_n, NET_143, VCC, SIM_RST);
    U74LVC07 U8028(NET_148, __A08_1___RL2_n, NET_145, __A08_1___Z2_n, NET_138, __A08_1___RL2_n, GND, __A08_1___RL2_n, NET_180, __A08_1___G2_n, NET_162, __A08_1___G2_n, NET_169, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U8029(NET_144, WZG_n, WL02_n, NET_145, NET_144, NET_146, GND, __A08_1___Z2_n, CZG, NET_146, RZG_n, __A08_1___Z2_n, NET_149, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U8030(NET_183, WBG_n, WL02_n, __A08_1___B2_n, NET_183, NET_184, GND, __A08_1___B2_n, CBG, NET_184, RBLG_n, __A08_1___B2_n, NET_182, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U8031(NET_182, NET_181, NET_168, NET_167, G02, NET_169, GND, NET_263, GND, XUY06_n, __A08_2___XUY2, NET_180, NET_161, VCC, SIM_RST);
    U74HC02 U8032(NET_181, NET_184, RCG_n, NET_164, WL01_n, WG3G_n, GND, WL03_n, WG4G_n, NET_163, L2GDG_n, L01_n, NET_168, VCC, SIM_RST);
    wire U8033_11_NC;
    wire U8033_12_NC;
    wire U8033_13_NC;
    U74HC02 U8033(NET_167, WG1G_n, WL02_n, G02, __A08_1___G2_n, CGG, GND, RGG_n, __A08_1___G2_n, NET_161, U8033_11_NC, U8033_12_NC, U8033_13_NC, VCC, SIM_RST);
    wire U8034_10_NC;
    wire U8034_11_NC;
    wire U8034_12_NC;
    wire U8034_13_NC;
    U74HC04 U8034(__A08_1___G2_n, __A08_1___GEM2, __A08_1___RL2_n, __A08_1___WL2, __A08_1___WL2, WL02_n, GND, __A08_1___MWL2, __A08_1___RL2_n, U8034_10_NC, U8034_11_NC, U8034_12_NC, U8034_13_NC, VCC, SIM_RST);
    U74HC02 U8035(NET_298, A2XG_n, __A08_2___A1_n, NET_294, WYLOG_n, WL03_n, GND, WL02_n, WYDG_n, NET_293, __A08_2__Y1_n, CUG, __A08_2__Y1, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U8036(MONEX, NET_298, __A08_2__X1_n, CLXC, CUG, __A08_2__X1, GND, __A08_2__Y1_n, NET_294, NET_293, __A08_2__Y1, __A08_2__X1_n, __A08_2__X1, VCC, SIM_RST);
    U74HC02 U8037(NET_302, __A08_2__X1_n, __A08_2__Y1_n, __A08_2___XUY1, __A08_2__X1, __A08_2__Y1, GND, NET_302, __A08_2___XUY1, NET_299, NET_302, __A08_2___SUMA1, __A08_2___CI_INTERNAL, VCC, SIM_RST);
    wire U8038_1_NC;
    wire U8038_2_NC;
    wire U8038_12_NC;
    wire U8038_13_NC;
    U74HC27 U8038(U8038_1_NC, U8038_2_NC, __A08_2___SUMA1, __A08_2___SUMB1, RULOG_n, NET_280, GND, NET_284, XUY05_n, __A08_2___XUY1, __A08_2___CI_IN, U8038_12_NC, U8038_13_NC, VCC, SIM_RST);
    U74HC04 U8039(__A08_2___CI_IN, NET_300, __A08_2___G1_n, __A08_2___GEM1, __A08_2___RL1_n, __A08_2___WL1, GND, WL03_n, __A08_2___WL1, __A08_2___MWL1, __A08_2___RL1_n, NET_250, __A08_2___CI_INTERNAL, VCC, SIM_RST);
    U74HC02 U8040(__A08_2___SUMB1, NET_299, NET_300, NET_283, WAG_n, WL03_n, GND, WL05_n, WALSG_n, NET_285, __A08_2___A1_n, CAG, NET_281, VCC, SIM_RST);
    U74LVC07 U8041(NET_284, CO06, NET_279, __A08_2___RL1_n, NET_291, __A08_2___L1_n, GND, __A08_2___Z1_n, NET_314, __A08_2___RL1_n, NET_315, __A08_2___RL1_n, NET_313, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U8042(NET_283, NET_285, NET_280, NET_278, CH03, NET_279, GND, NET_291, NET_282, NET_289, NET_290, __A08_2___A1_n, NET_281, VCC, SIM_RST);
    U74HC02 U8043(NET_278, RAG_n, __A08_2___A1_n, NET_282, WLG_n, WL03_n, GND, G06_n, G2LSG_n, NET_289, __A08_2___L1_n, CLG1G, NET_290, VCC, SIM_RST);
    wire U8044_1_NC;
    wire U8044_2_NC;
    wire U8044_3_NC;
    wire U8044_4_NC;
    wire U8044_5_NC;
    wire U8044_6_NC;
    wire U8044_12_NC;
    wire U8044_13_NC;
    U74HC27 U8044(U8044_1_NC, U8044_2_NC, U8044_3_NC, U8044_4_NC, U8044_5_NC, U8044_6_NC, GND, __A08_2___RL_OUT_1, RLG_n, __A08_2___L1_n, GND, U8044_12_NC, U8044_13_NC, VCC, SIM_RST);
    wire U8045_1_NC;
    wire U8045_2_NC;
    wire U8045_3_NC;
    U74HC02 #(0, 0, 1, 0) U8045(U8045_1_NC, U8045_2_NC, U8045_3_NC, NET_287, WQG_n, WL03_n, GND, NET_287, NET_286, __A08_2___Q1_n, __A08_2___Q1_n, CQG, NET_286, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U8046(NET_288, RQG_n, __A08_2___Q1_n, NET_317, WZG_n, WL03_n, GND, NET_317, NET_316, NET_314, __A08_2___Z1_n, CZG, NET_316, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U8047(NET_312, RZG_n, __A08_2___Z1_n, NET_321, WBG_n, WL03_n, GND, NET_321, NET_322, __A08_2___B1_n, __A08_2___B1_n, CBG, NET_322, VCC, SIM_RST);
    U74HC02 U8048(NET_319, RBLG_n, __A08_2___B1_n, NET_320, NET_322, RCG_n, GND, WL02_n, WG3G_n, NET_309, WL04_n, WG4G_n, NET_308, VCC, SIM_RST);
    U74HC27 U8049(__A08_2___RL_OUT_1, NET_288, MDT03, R1C, R15, NET_313, GND, NET_318, NET_319, NET_320, NET_305, NET_315, NET_312, VCC, SIM_RST);
    U74LVC07 U8050(NET_263, CO06, NET_318, __A08_2___RL1_n, NET_304, __A08_2___G1_n, GND, __A08_2___G1_n, NET_303, __A08_2___RL2_n, NET_230, L04_n, NET_240, VCC, SIM_RST);
    U74HC02 U8051(NET_307, L2GDG_n, L02_n, NET_306, WG1G_n, WL03_n, GND, __A08_2___G1_n, CGG, G03, RGG_n, __A08_2___G1_n, NET_305, VCC, SIM_RST);
    U74HC4002 #(1, 0) U8052(NET_304, G03ED, SA03, NET_309, NET_308, NET_311, GND, NET_310, G04ED, SA04, NET_257, NET_256, NET_255, VCC, SIM_RST);
    wire U8053_3_NC;
    wire U8053_4_NC;
    wire U8053_5_NC;
    wire U8053_6_NC;
    wire U8053_8_NC;
    wire U8053_9_NC;
    wire U8053_10_NC;
    wire U8053_11_NC;
    U74HC27 #(1, 0, 0) U8053(NET_307, NET_306, U8053_3_NC, U8053_4_NC, U8053_5_NC, U8053_6_NC, GND, U8053_8_NC, U8053_9_NC, U8053_10_NC, U8053_11_NC, NET_303, G03, VCC, SIM_RST);
    U74HC02 U8054(NET_251, A2XG_n, __A08_2___A2_n, NET_253, WYLOG_n, WL04_n, GND, WL03_n, WYDG_n, NET_252, __A08_2__Y2_n, CUG, __A08_2__Y2, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U8055(MONEX, NET_251, __A08_2__X2_n, CLXC, CUG, __A08_2__X2, GND, __A08_2__Y2_n, NET_253, NET_252, __A08_2__Y2, __A08_2__X2_n, __A08_2__X2, VCC, SIM_RST);
    wire U8056_8_NC;
    wire U8056_9_NC;
    wire U8056_10_NC;
    U74HC02 U8056(NET_245, __A08_2__X2_n, __A08_2__Y2_n, __A08_2___XUY2, __A08_2__X2, __A08_2__Y2, GND, U8056_8_NC, U8056_9_NC, U8056_10_NC, NET_245, __A08_2___XUY2, NET_248, VCC, SIM_RST);
    wire U8057_1_NC;
    wire U8057_2_NC;
    wire U8057_12_NC;
    wire U8057_13_NC;
    U74HC27 U8057(U8057_1_NC, U8057_2_NC, NET_245, __A08_2___SUMA2, __A08_2___CO_IN, CI05_n, GND, NET_249, __A08_2___SUMA2, __A08_2___SUMB2, RULOG_n, U8057_12_NC, U8057_13_NC, VCC, SIM_RST);
    U74HC02 U8058(__A08_2___SUMB2, NET_248, NET_250, NET_234, WAG_n, WL04_n, GND, WL06_n, WALSG_n, NET_233, __A08_2___A2_n, CAG, NET_232, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U8059(NET_234, NET_233, NET_249, NET_235, CH04, NET_230, GND, NET_240, NET_268, NET_269, NET_270, __A08_2___A2_n, NET_232, VCC, SIM_RST);
    U74HC02 U8060(NET_235, RAG_n, __A08_2___A2_n, NET_268, WLG_n, WL04_n, GND, G07_n, G2LSG_n, NET_269, L04_n, CLG1G, NET_270, VCC, SIM_RST);
    U74HC27 U8061(RLG_n, L04_n, __A08_2___RL_OUT_2, NET_236, NET_242, NET_241, GND, NET_231, MDT04, R1C, R15, __A08_2___RL_OUT_2, GND, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U8062(NET_272, WQG_n, WL04_n, __A08_2___Q2_n, NET_272, NET_271, GND, __A08_2___Q2_n, CQG, NET_271, RQG_n, __A08_2___Q2_n, NET_236, VCC, SIM_RST);
    U74LVC07 U8063(NET_241, __A08_2___RL2_n, NET_238, __A08_2___Z2_n, NET_231, __A08_2___RL2_n, GND, __A08_2___RL2_n, NET_273, __A08_2___G2_n, NET_255, __A08_2___G2_n, NET_262, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U8064(NET_237, WZG_n, WL04_n, NET_238, NET_237, NET_239, GND, __A08_2___Z2_n, CZG, NET_239, RZG_n, __A08_2___Z2_n, NET_242, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U8065(NET_276, WBG_n, WL04_n, __A08_2___B2_n, NET_276, NET_277, GND, __A08_2___B2_n, CBG, NET_277, RBLG_n, __A08_2___B2_n, NET_275, VCC, SIM_RST);
    wire U8066_8_NC;
    wire U8066_9_NC;
    wire U8066_10_NC;
    wire U8066_11_NC;
    U74HC27 #(0, 1, 0) U8066(NET_275, NET_274, NET_261, NET_260, G04, NET_262, GND, U8066_8_NC, U8066_9_NC, U8066_10_NC, U8066_11_NC, NET_273, NET_254, VCC, SIM_RST);
    U74HC02 U8067(NET_274, NET_277, RCG_n, NET_257, WL03_n, WG3G_n, GND, WL05_n, WG4G_n, NET_256, L2GDG_n, __A08_2___L1_n, NET_261, VCC, SIM_RST);
    wire U8068_11_NC;
    wire U8068_12_NC;
    wire U8068_13_NC;
    U74HC02 U8068(NET_260, WG1G_n, WL04_n, G04, __A08_2___G2_n, CGG, GND, RGG_n, __A08_2___G2_n, NET_254, U8068_11_NC, U8068_12_NC, U8068_13_NC, VCC, SIM_RST);
    wire U8069_10_NC;
    wire U8069_11_NC;
    wire U8069_12_NC;
    wire U8069_13_NC;
    U74HC04 U8069(__A08_2___G2_n, __A08_2___GEM2, __A08_2___RL2_n, __A08_2___WL2, __A08_2___WL2, WL04_n, GND, __A08_2___MWL2, __A08_2___RL2_n, U8069_10_NC, U8069_11_NC, U8069_12_NC, U8069_13_NC, VCC, SIM_RST);
    U74HC4002 U8070(__A08_1___SUMA1, NET_209, XUY01_n, CI01_n, GND, NET_174, GND, NET_173, NET_152, XUY02_n, __A08_1___CI_INTERNAL, WHOMP, __A08_1___SUMA2, VCC, SIM_RST);
    U74HC4002 U8071(__A08_2___SUMA1, NET_302, __A08_2___XUY1, __A08_2___CI_IN, GND, NET_267, GND, NET_266, NET_245, __A08_2___XUY2, __A08_2___CI_INTERNAL, WHOMP, __A08_2___SUMA2, VCC, SIM_RST);
endmodule