`include "components/agc_parts.v"

module timer(VCC, GND, SIM_RST, CLOCK, STOP, PHS2, PHS2_n, PHS3_n, PHS4, PHS4_n, RT, RT_n, WT, WT_n, CT, CT_n, TT_n, OVFSTB_n, CLK, P01, P01_n, P02, P02_n, P03, P03_n, P04, P04_n, P05, P05_n);
    input wire SIM_RST;
    output wire RT;
    wire __A02_1__cdiv_1__B;
    wire __A02_1__cdiv_2__F;
    wire NET_61;
    output wire PHS4;
    input wire VCC;
    wire __A02_2__F01D;
    wire __A02_1__oddset;
    wire __A02_1__ovfstb_r4;
    output wire P01_n;
    output wire P05_n;
    wire __A02_1__cdiv_1__D;
    wire __A02_1__ovfstb_r3;
    output wire PHS2;
    output wire P05;
    output wire P04_n;
    wire __A02_1__RINGB_n;
    wire __A02_1__evnset;
    output wire P04;
    wire NET_43;
    wire NET_58;
    wire NET_57;
    wire __A02_1__cdiv_2__FS;
    wire __A02_1__cdiv_2__C;
    wire __A02_1__ovfstb_r1;
    wire NET_62;
    output wire PHS3_n;
    output wire CT_n;
    wire __A02_2__F01C;
    wire __A02_1__cdiv_2__FS_n;
    input wire STOP;
    output wire P01;
    wire __A02_1__Q2A;
    wire NET_56;
    wire NET_65;
    wire __A02_2__F01A;
    wire __A02_1__cdiv_1__FS_n;
    output wire CLK;
    output wire P03_n;
    wire __A02_1__ovfstb_r6;
    wire __A02_1__ovfstb_r2;
    wire __A02_1__cdiv_1__A;
    wire __A02_1__cdiv_1__FS;
    wire __A02_1__ovfstb_r5;
    output wire P03;
    wire __A02_1__MONWT;
    output wire P02_n;
    wire NET_63;
    wire __A02_1__cdiv_2__D;
    output wire PHS2_n;
    wire NET_64;
    output wire TT_n;
    output wire WT;
    output wire RT_n;
    wire NET_60;
    wire NET_59;
    wire __A02_1__cdiv_2__B;
    wire __A02_1__cdiv_2__A;
    wire __A02_2__FS01;
    output wire PHS4_n;
    output wire CT;
    wire __A02_1__EVNSET_n;
    input wire GND;
    wire __A02_1__ODDSET_n;
    wire __A02_2__F01B;
    wire __A02_1__RINGA_n;
    output wire WT_n;
    output wire OVFSTB_n;
    input wire CLOCK;
    wire __A02_2__FS01_n;
    output wire P02;

    U74HC02 #(0, 1, 0, 0) U12(P01, NET_57, P01_n, P01_n, P01, NET_56, GND, __A02_1__RINGA_n, P01, NET_65, P01_n, __A02_1__RINGB_n, NET_63, VCC, SIM_RST);
    U74HC04 U5(__A02_1__cdiv_1__FS_n, WT, WT, WT_n, WT, TT_n, GND, __A02_1__ovfstb_r5, __A02_1__ovfstb_r4, __A02_1__ovfstb_r6, __A02_1__ovfstb_r5, OVFSTB_n, __A02_1__ovfstb_r2, VCC, SIM_RST);
    wire U2_8_NC;
    wire U2_9_NC;
    wire U2_10_NC;
    wire U2_11_NC;
    U74HC27 #(0, 1, 0) U2(__A02_1__cdiv_1__D, CLOCK, __A02_1__cdiv_1__B, CLOCK, PHS2, __A02_1__cdiv_1__A, GND, U2_8_NC, U2_9_NC, U2_10_NC, U2_11_NC, __A02_1__cdiv_1__B, __A02_1__cdiv_1__A, VCC, SIM_RST);
    wire U10_12_NC;
    wire U10_13_NC;
    U74HC04 U10(CT, PHS3_n, WT_n, CLK, WT_n, __A02_1__MONWT, GND, __A02_1__Q2A, WT_n, RT_n, RT, U10_12_NC, U10_13_NC, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U17(__A02_2__F01D, __A02_2__FS01_n, __A02_2__F01B, __A02_2__FS01_n, __A02_2__F01B, __A02_2__FS01, GND, __A02_2__FS01_n, __A02_2__F01A, __A02_2__FS01, __A02_2__F01A, __A02_2__FS01, __A02_2__F01C, VCC, SIM_RST);
    U74HC02 U9(__A02_1__ovfstb_r1, CT_n, __A02_1__ovfstb_r2, __A02_1__ovfstb_r2, __A02_1__ovfstb_r6, __A02_1__ovfstb_r1, GND, __A02_1__ovfstb_r4, __A02_1__ovfstb_r2, __A02_1__ovfstb_r3, __A02_1__ovfstb_r3, __A02_1__ovfstb_r1, __A02_1__ovfstb_r4, VCC, SIM_RST);
    wire U18_8_NC;
    wire U18_9_NC;
    wire U18_10_NC;
    wire U18_11_NC;
    U74HC27 #(0, 1, 0) U18(__A02_2__F01D, P01_n, __A02_2__F01B, P01_n, __A02_2__F01C, __A02_2__F01A, GND, U18_8_NC, U18_9_NC, U18_10_NC, U18_11_NC, __A02_2__F01B, __A02_2__F01A, VCC, SIM_RST);
    wire U11_8_NC;
    wire U11_9_NC;
    wire U11_10_NC;
    wire U11_11_NC;
    U74HC27 U11(__A02_1__RINGB_n, P05_n, P04, P05, __A02_1__RINGA_n, NET_56, GND, U11_8_NC, U11_9_NC, U11_10_NC, U11_11_NC, NET_57, P04_n, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U15(P04, NET_60, P04_n, P04_n, P04, NET_62, GND, __A02_1__RINGB_n, P04, NET_59, P04_n, __A02_1__RINGA_n, NET_58, VCC, SIM_RST);
    U74HC04 U3(__A02_1__cdiv_1__D, __A02_1__cdiv_2__F, PHS2, PHS2_n, PHS4, PHS4_n, GND, NET_43, __A02_1__cdiv_1__B, CT, NET_43, CT_n, CT, VCC, SIM_RST);
    U74HC04 U8(__A02_1__cdiv_2__D, __A02_1__RINGA_n, __A02_1__oddset, __A02_1__ODDSET_n, __A02_1__cdiv_2__C, __A02_1__RINGB_n, GND, __A02_1__evnset, __A02_1__RINGB_n, __A02_1__EVNSET_n, __A02_1__evnset, RT, __A02_1__cdiv_1__A, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U14(P03, NET_61, P03_n, P03_n, P03, NET_64, GND, __A02_1__RINGA_n, P03, NET_60, P03_n, __A02_1__RINGB_n, NET_62, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U1(__A02_1__cdiv_1__D, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__B, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__B, __A02_1__cdiv_1__FS, GND, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__A, __A02_1__cdiv_1__FS, __A02_1__cdiv_1__A, __A02_1__cdiv_1__FS, PHS2, VCC, SIM_RST);
    wire U7_8_NC;
    wire U7_9_NC;
    wire U7_10_NC;
    wire U7_11_NC;
    U74HC27 #(0, 1, 0) U7(__A02_1__cdiv_2__D, __A02_1__cdiv_2__F, __A02_1__cdiv_2__B, __A02_1__cdiv_2__F, __A02_1__cdiv_2__C, __A02_1__cdiv_2__A, GND, U7_8_NC, U7_9_NC, U7_10_NC, U7_11_NC, __A02_1__cdiv_2__B, __A02_1__cdiv_2__A, VCC, SIM_RST);
    wire U16_8_NC;
    wire U16_9_NC;
    wire U16_10_NC;
    wire U16_11_NC;
    wire U16_12_NC;
    wire U16_13_NC;
    U74HC02 #(0, 1, 0, 0) U16(P05, NET_59, P05_n, P05_n, P05, NET_58, GND, U16_8_NC, U16_9_NC, U16_10_NC, U16_11_NC, U16_12_NC, U16_13_NC, VCC, SIM_RST);
    wire U4_8_NC;
    wire U4_9_NC;
    wire U4_10_NC;
    wire U4_11_NC;
    wire U4_12_NC;
    wire U4_13_NC;
    U74HC02 U4(PHS4, __A02_1__cdiv_2__F, __A02_1__cdiv_1__A, __A02_1__oddset, STOP, __A02_1__RINGA_n, GND, U4_8_NC, U4_9_NC, U4_10_NC, U4_11_NC, U4_12_NC, U4_13_NC, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U6(__A02_1__cdiv_2__D, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__FS, GND, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__A, __A02_1__cdiv_2__FS, __A02_1__cdiv_2__A, __A02_1__cdiv_2__FS, __A02_1__cdiv_2__C, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U13(P02, NET_65, P02_n, P02_n, P02, NET_63, GND, __A02_1__RINGB_n, P02, NET_61, P02_n, __A02_1__RINGA_n, NET_64, VCC, SIM_RST);
endmodule