`timescale 1ns/1ps
`default_nettype none

module rupt_service(SIM_RST, SIM_CLK, p4VSW, GND, GOJAM, T10, S10, S10_n, S11_n, S12_n, WL01_n, WL02_n, WL03_n, WL09_n, WL10_n, WL11_n, WL12_n, WL13_n, WL14_n, WL16_n, SUMA01_n, SUMB01_n, SUMA02_n, SUMB02_n, SUMA03_n, SUMB03_n, SUMA11_n, SUMB11_n, SUMA12_n, SUMB12_n, SUMA13_n, SUMB13_n, SUMA14_n, SUMB14_n, SUMA16_n, SUMB16_n, XB0_n, XB1_n, XB4_n, XB6_n, XB7_n, XT0_n, XT1_n, XT2_n, XT3_n, XT4_n, XT5_n, E5, E6, E7_n, STRGAT, CEBG, CFBG, OVF_n, R6, RB1F, RBBEG_n, REBG_n, RFBG_n, RRPA, RSTRT, U2BBKG_n, WBBEG_n, WEBG_n, WFBG_n, WOVR_n, ZOUT_n, DLKPLS, HNDRPT, KRPT, KYRPT1, KYRPT2, RADRPT, UPRUPT, CA2_n, CA3_n, CAD1, CAD2, CAD3, CAD4, CAD5, CAD6, MKRPT, EB9, EB10, EB11_n, RL01_n, RL02_n, RL03_n, RL04_n, RL05_n, RL06_n, RL09_n, RL10_n, RL11_n, RL12_n, RL13_n, RL14_n, RL15_n, RL16_n, RUPTOR_n, ROPER, ROPES, ROPET, HIMOD, LOMOD, STR19, STR210, STR311, STR412, STR14, STR58, STR912, T6RPT, DRPRST);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VSW;
    input wire GND;
    input wire CA2_n;
    input wire CA3_n;
    input wire CAD1;
    input wire CAD2;
    input wire CAD3;
    input wire CAD4;
    input wire CAD5;
    input wire CAD6;
    input wire CEBG;
    input wire CFBG;
    input wire DLKPLS;
    output wire DRPRST;
    input wire E5;
    input wire E6;
    input wire E7_n;
    output wire EB10;
    output wire EB11_n;
    output wire EB9;
    input wire GOJAM;
    output wire HIMOD;
    input wire HNDRPT;
    input wire KRPT;
    input wire KYRPT1;
    input wire KYRPT2;
    output wire LOMOD;
    input wire MKRPT;
    input wire OVF_n;
    input wire R6;
    input wire RADRPT;
    input wire RB1F;
    input wire RBBEG_n;
    input wire REBG_n;
    input wire RFBG_n;
    output wire RL01_n; //FPGA#wand
    output wire RL02_n; //FPGA#wand
    output wire RL03_n; //FPGA#wand
    output wire RL04_n; //FPGA#wand
    output wire RL05_n; //FPGA#wand
    output wire RL06_n; //FPGA#wand
    output wire RL09_n; //FPGA#wand
    output wire RL10_n; //FPGA#wand
    output wire RL11_n; //FPGA#wand
    output wire RL12_n; //FPGA#wand
    output wire RL13_n; //FPGA#wand
    output wire RL14_n; //FPGA#wand
    output wire RL15_n; //FPGA#wand
    output wire RL16_n; //FPGA#wand
    output wire ROPER;
    output wire ROPES;
    output wire ROPET;
    input wire RRPA;
    input wire RSTRT;
    output wire RUPTOR_n;
    input wire S10;
    input wire S10_n;
    input wire S11_n;
    input wire S12_n;
    output wire STR14;
    output wire STR19;
    output wire STR210;
    output wire STR311;
    output wire STR412;
    output wire STR58;
    output wire STR912;
    input wire STRGAT;
    input wire SUMA01_n;
    input wire SUMA02_n;
    input wire SUMA03_n;
    input wire SUMA11_n;
    input wire SUMA12_n;
    input wire SUMA13_n;
    input wire SUMA14_n;
    input wire SUMA16_n;
    input wire SUMB01_n;
    input wire SUMB02_n;
    input wire SUMB03_n;
    input wire SUMB11_n;
    input wire SUMB12_n;
    input wire SUMB13_n;
    input wire SUMB14_n;
    input wire SUMB16_n;
    input wire T10;
    output wire T6RPT;
    input wire U2BBKG_n;
    input wire UPRUPT;
    input wire WBBEG_n;
    input wire WEBG_n;
    input wire WFBG_n;
    input wire WL01_n;
    input wire WL02_n;
    input wire WL03_n;
    input wire WL09_n;
    input wire WL10_n;
    input wire WL11_n;
    input wire WL12_n;
    input wire WL13_n;
    input wire WL14_n;
    input wire WL16_n;
    input wire WOVR_n;
    input wire XB0_n;
    input wire XB1_n;
    input wire XB4_n;
    input wire XB6_n;
    input wire XB7_n;
    input wire XT0_n;
    input wire XT1_n;
    input wire XT2_n;
    input wire XT3_n;
    input wire XT4_n;
    input wire XT5_n;
    input wire ZOUT_n;
    wire __A15_1__BBK1;
    wire __A15_1__BBK2;
    wire __A15_1__BBK3;
    wire __A15_1__BK16;
    wire __A15_1__DNRPTA;
    wire __A15_1__EB10_n;
    wire __A15_1__EB11;
    wire __A15_1__EB9_n;
    wire __A15_1__F11;
    wire __A15_1__F11_n;
    wire __A15_1__F12;
    wire __A15_1__F12_n;
    wire __A15_1__F13;
    wire __A15_1__F13_n;
    wire __A15_1__F14;
    wire __A15_1__F14_n;
    wire __A15_1__F15;
    wire __A15_1__F15_n;
    wire __A15_1__F16;
    wire __A15_1__F16_n;
    wire __A15_1__FB11;
    wire __A15_1__FB11_n;
    wire __A15_1__FB12;
    wire __A15_1__FB12_n;
    wire __A15_1__FB13;
    wire __A15_1__FB13_n;
    wire __A15_1__FB14;
    wire __A15_1__FB14_n;
    wire __A15_1__FB16;
    wire __A15_1__FB16_n;
    wire __A15_1__KRPTA_n;
    wire __A15_1__PRPOR1;
    wire __A15_1__PRPOR2;
    wire __A15_1__PRPOR3;
    wire __A15_1__PRPOR4;
    wire __A15_1__RPTA12;
    wire __A15_1__RPTAD6;
    wire __A15_1__RRPA1_n;
    wire __A15_2__036H;
    wire __A15_2__036L;
    wire __A15_2__147H;
    wire __A15_2__147L;
    wire __A15_2__2510H;
    wire __A15_2__2510L;
    wire __A15_2__KY1RST;
    wire __A15_2__KY2RST;
    wire __A15_2__NE00;
    wire __A15_2__NE01;
    wire __A15_2__NE012_n;
    wire __A15_2__NE02;
    wire __A15_2__NE03;
    wire __A15_2__NE036_n;
    wire __A15_2__NE04;
    wire __A15_2__NE05;
    wire __A15_2__NE06;
    wire __A15_2__NE07;
    wire __A15_2__NE10;
    wire __A15_2__NE147_n;
    wire __A15_2__NE2510_n;
    wire __A15_2__NE345_n;
    wire __A15_2__NE6710_n;
    wire __A15_2__RPTAD3;
    wire __A15_2__RPTAD4;
    wire __A15_2__RPTAD5;
    wire __A15_NET_149;
    wire __A15_NET_150;
    wire __A15_NET_151;
    wire __A15_NET_152;
    wire __A15_NET_153;
    wire __A15_NET_154;
    wire __A15_NET_155;
    wire __A15_NET_156;
    wire __A15_NET_157;
    wire __A15_NET_158;
    wire __A15_NET_159;
    wire __A15_NET_160;
    wire __A15_NET_161;
    wire __A15_NET_162;
    wire __A15_NET_163;
    wire __A15_NET_164;
    wire __A15_NET_165;
    wire __A15_NET_166;
    wire __A15_NET_167;
    wire __A15_NET_168;
    wire __A15_NET_171;
    wire __A15_NET_174;
    wire __A15_NET_175;
    wire __A15_NET_176;
    wire __A15_NET_177;
    wire __A15_NET_179;
    wire __A15_NET_181;
    wire __A15_NET_184;
    wire __A15_NET_185;
    wire __A15_NET_186;
    wire __A15_NET_187;
    wire __A15_NET_188;
    wire __A15_NET_189;
    wire __A15_NET_192;
    wire __A15_NET_195;
    wire __A15_NET_197;
    wire __A15_NET_198;
    wire __A15_NET_199;
    wire __A15_NET_200;
    wire __A15_NET_201;
    wire __A15_NET_202;
    wire __A15_NET_203;
    wire __A15_NET_204;
    wire __A15_NET_205;
    wire __A15_NET_206;
    wire __A15_NET_207;
    wire __A15_NET_208;
    wire __A15_NET_209;
    wire __A15_NET_210;
    wire __A15_NET_213;
    wire __A15_NET_214;
    wire __A15_NET_215;
    wire __A15_NET_216;
    wire __A15_NET_217;
    wire __A15_NET_218;
    wire __A15_NET_219;
    wire __A15_NET_220;
    wire __A15_NET_221;
    wire __A15_NET_222;
    wire __A15_NET_223;
    wire __A15_NET_224;
    wire __A15_NET_225;
    wire __A15_NET_226;
    wire __A15_NET_227;
    wire __A15_NET_228;
    wire __A15_NET_229; //FPGA#wand
    wire __A15_NET_232; //FPGA#wand
    wire __A15_NET_234;
    wire __A15_NET_235;
    wire __A15_NET_236;
    wire __A15_NET_237;
    wire __A15_NET_238;
    wire __A15_NET_239;
    wire __A15_NET_240;
    wire __A15_NET_241;
    wire __A15_NET_242;
    wire __A15_NET_243;
    wire __A15_NET_244;
    wire __A15_NET_245;
    wire __A15_NET_246;
    wire __A15_NET_251;
    wire __A15_NET_260;
    wire __A15_NET_261;
    wire __A15_NET_262;
    wire __A15_NET_265;
    wire __A15_NET_266;
    wire __A15_NET_267;
    wire __A15_NET_268;
    wire __A15_NET_269;
    wire __A15_NET_270;
    wire __A15_NET_271;
    wire __A15_NET_272;
    wire __A15_NET_273;
    wire __A15_NET_274;
    wire __A15_NET_282;
    wire __A15_NET_283;
    wire __A15_NET_284;
    wire __A15_NET_285;
    wire __A15_NET_286;
    wire __A15_NET_287;
    wire __A15_NET_290;
    wire __A15_NET_291;
    wire __A15_NET_294;
    wire __A15_NET_295;
    wire __A15_NET_296;
    wire __A15_NET_297;
    wire __A15_NET_298;
    wire __A15_NET_299;
    wire __A15_NET_300;
    wire __A15_NET_301;
    wire __A15_NET_302;
    wire __A15_NET_303;
    wire __A15_NET_304;
    wire __A15_NET_305;
    wire __A15_NET_306;
    wire __A15_NET_307;
    wire __A15_NET_310;

    pullup R15001(__A15_NET_229);
    pullup R15002(__A15_NET_232);
    U74HC02 U15001(__A15_NET_200, WL16_n, WFBG_n, __A15_1__FB16, __A15_1__FB16_n, CFBG, GND, __A15_1__FB16_n, RFBG_n, __A15_1__BK16, WL14_n, WFBG_n, __A15_NET_198, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0, 1'b0) U15002(__A15_NET_200, __A15_NET_201, SUMA16_n, U2BBKG_n, SUMB16_n, __A15_NET_201, GND, __A15_NET_199, SUMA14_n, U2BBKG_n, SUMB14_n, __A15_1__FB16_n, __A15_1__FB16, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15003(__A15_1__BK16, __A15_NET_195, __A15_1__BK16, __A15_NET_197, __A15_NET_206, __A15_NET_207, GND, __A15_NET_202, __A15_NET_204, __A15_NET_192, __A15_NET_165, __A15_NET_210, __A15_NET_149, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U15004(__A15_NET_195, RL16_n, __A15_NET_197, RL15_n, __A15_NET_207, RL14_n, GND, RL13_n, __A15_NET_202, RL12_n, __A15_NET_189, RL11_n, __A15_NET_188, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 #(1'b1, 1'b0, 1'b1, 1'b0) U15005(__A15_NET_198, __A15_NET_199, SUMA13_n, U2BBKG_n, SUMB13_n, __A15_NET_209, GND, __A15_1__FB13_n, __A15_NET_208, __A15_NET_209, __A15_1__FB13, __A15_1__FB14_n, __A15_1__FB14, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15006(__A15_1__FB14, __A15_1__FB14_n, CFBG, __A15_NET_206, __A15_1__FB14_n, RFBG_n, GND, WL13_n, WFBG_n, __A15_NET_208, __A15_1__FB13_n, CFBG, __A15_1__FB13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15007(__A15_NET_204, __A15_1__FB13_n, RFBG_n, __A15_NET_203, WL12_n, WFBG_n, GND, __A15_1__FB12_n, CFBG, __A15_1__FB12, __A15_1__FB12_n, RFBG_n, __A15_NET_161, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0, 1'b0) U15008(SUMA12_n, U2BBKG_n, __A15_NET_203, __A15_NET_205, __A15_1__FB12, __A15_1__FB12_n, GND, __A15_NET_189, RSTRT, __A15_NET_161, __A15_1__RPTA12, __A15_NET_205, SUMB12_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15009(__A15_NET_162, WFBG_n, WL11_n, __A15_1__FB11, __A15_1__FB11_n, CFBG, GND, __A15_1__FB11_n, RFBG_n, __A15_NET_157, __A15_NET_157, __A15_NET_166, __A15_NET_188, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0, 1'b0) U15010(SUMA11_n, U2BBKG_n, __A15_NET_162, __A15_NET_163, __A15_1__FB11, __A15_1__FB11_n, GND, __A15_NET_158, SUMA03_n, U2BBKG_n, SUMB03_n, __A15_NET_163, SUMB11_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15011(__A15_NET_159, WL11_n, WEBG_n, __A15_NET_160, WL03_n, WBBEG_n, GND, EB11_n, CEBG, __A15_1__EB11, REBG_n, EB11_n, __A15_NET_166, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1, 1'b0) U15012(EB11_n, __A15_NET_158, __A15_NET_159, __A15_NET_160, __A15_1__EB11,  , GND,  , __A15_NET_167, __A15_NET_168, __A15_NET_164, EB10, __A15_1__EB10_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15013(__A15_1__BBK3, EB11_n, RBBEG_n, __A15_NET_168, WL10_n, WEBG_n, GND, WL02_n, WBBEG_n, __A15_NET_164, __A15_1__EB10_n, CEBG, EB10, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15014(SUMA02_n, U2BBKG_n, SUMA01_n, U2BBKG_n, SUMB01_n, __A15_NET_150, GND, __A15_1__F14, __A15_NET_153, __A15_NET_154, __A15_1__FB14_n, __A15_NET_167, SUMB02_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15015(__A15_NET_165, REBG_n, __A15_1__EB10_n, __A15_1__BBK2, __A15_1__EB10_n, RBBEG_n, GND, WL09_n, WEBG_n, __A15_NET_151, WL01_n, WBBEG_n, __A15_NET_152, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U15016(__A15_NET_192, RL10_n, __A15_NET_210, RL09_n, __A15_NET_181, RL06_n, GND, __A15_NET_229, __A15_NET_294, __A15_NET_229, __A15_NET_296, __A15_NET_232, __A15_NET_291, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC4002 #(1'b1, 1'b1, 1'b0) U15017(__A15_1__EB9_n, __A15_NET_150, __A15_NET_151, __A15_NET_152, EB9,  , GND,  , __A15_1__FB14_n, __A15_1__FB16_n, E7_n, __A15_NET_153, __A15_1__F16, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15018(EB9, __A15_1__EB9_n, CEBG, __A15_NET_149, REBG_n, __A15_1__EB9_n, GND, __A15_1__EB9_n, RBBEG_n, __A15_1__BBK1, __A15_1__FB11_n, __A15_NET_153, __A15_NET_155, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15019(S12_n, __A15_NET_153, __A15_1__F11_n, __A15_1__F11, __A15_1__F12_n, __A15_1__F12, GND, __A15_1__F13_n, __A15_1__F13, __A15_1__F14_n, __A15_1__F14, __A15_1__F15_n, __A15_1__F15, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15020(__A15_1__F11_n, __A15_NET_155, __A15_NET_156, __A15_NET_156, S11_n, S12_n, GND, __A15_NET_153, __A15_1__FB12, __A15_1__F12_n, __A15_NET_153, __A15_1__FB13_n, __A15_1__F13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15021(E5, __A15_1__FB16_n, __A15_1__FB16_n, __A15_NET_184, __A15_NET_153, __A15_1__F15, GND, __A15_NET_184, E7_n, __A15_1__FB14_n, E6, __A15_NET_154, E7_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15022(__A15_1__F16, __A15_1__F16_n, __A15_NET_305, __A15_NET_301, KRPT, __A15_1__KRPTA_n, GND, __A15_NET_245, __A15_NET_244, __A15_NET_213, __A15_NET_224, __A15_1__PRPOR1, __A15_NET_218, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15023(XB4_n, XT4_n, __A15_1__KRPTA_n, XB0_n, XT5_n, __A15_NET_186, GND, __A15_NET_175, __A15_NET_185, __A15_NET_187, GOJAM, __A15_NET_187, __A15_1__KRPTA_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b0, 1'b0) U15024(__A15_NET_185, RADRPT, __A15_NET_175, __A15_NET_174, HNDRPT, __A15_NET_171, GND, __A15_NET_179, __A15_1__RRPA1_n, __A15_1__RPTAD6, __A15_1__RRPA1_n, __A15_NET_177, __A15_1__RPTA12, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15025(__A15_NET_174, __A15_NET_186, __A15_1__PRPOR1, __A15_NET_185, __A15_1__DNRPTA, __A15_1__PRPOR3, GND, __A15_NET_179, __A15_1__PRPOR2, __A15_1__PRPOR3, __A15_1__PRPOR4, __A15_NET_171, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U15026(__A15_1__PRPOR4, __A15_1__PRPOR1, __A15_1__DNRPTA, __A15_NET_175, __A15_NET_174,  , GND,  , __A15_NET_171, __A15_NET_175, __A15_1__PRPOR1, __A15_1__DNRPTA, __A15_NET_177, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U15027(__A15_NET_181, CAD6, __A15_1__RPTAD6, __A15_NET_176, __A15_NET_177, RUPTOR_n, GND, __A15_NET_176, T10, RUPTOR_n, WOVR_n, OVF_n, __A15_NET_305, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15028(CA3_n, XB1_n, __A15_NET_306, GOJAM, __A15_NET_307, __A15_NET_295, GND, __A15_NET_307, XT0_n, XB4_n, __A15_1__KRPTA_n, T6RPT, ZOUT_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b1, 1'b0) U15029(__A15_NET_306, T6RPT, __A15_NET_295, __A15_NET_238, __A15_NET_302, __A15_NET_240, GND, __A15_NET_303, __A15_NET_243, __A15_NET_239, __A15_NET_236, __A15_NET_223, __A15_NET_237, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15030(CA3_n, XB0_n, __A15_NET_238, GOJAM, __A15_NET_300, __A15_NET_240, GND, __A15_NET_300, XB0_n, XT1_n, __A15_1__KRPTA_n, __A15_NET_302, __A15_NET_301, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15031(CA2_n, XB6_n, __A15_NET_239, GOJAM, __A15_NET_304, __A15_NET_243, GND, __A15_NET_304, XT1_n, XB4_n, __A15_1__KRPTA_n, __A15_NET_303, __A15_NET_301, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15032(CA2_n, XB7_n, __A15_NET_237, GOJAM, __A15_NET_235, __A15_NET_223, GND, __A15_NET_235, XT2_n, XB0_n, __A15_1__KRPTA_n, __A15_NET_236, __A15_NET_301, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b0, 1'b0) U15033(__A15_NET_234, KYRPT1, __A15_NET_225, __A15_NET_215, UPRUPT, __A15_NET_219, GND, DLKPLS, __A15_1__DNRPTA, __A15_NET_220, __A15_NET_295, __A15_NET_238, __A15_NET_241, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1, 1'b0) U15034(__A15_NET_234, GOJAM, XB4_n, XT2_n, __A15_1__KRPTA_n, __A15_2__KY1RST, GND, __A15_NET_226, KYRPT2, MKRPT, __A15_NET_217, __A15_NET_225, __A15_2__KY1RST, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15035(__A15_NET_226, GOJAM, XT3_n, XB0_n, __A15_1__KRPTA_n, __A15_2__KY2RST, GND, __A15_NET_219, __A15_NET_215, GOJAM, __A15_NET_246, __A15_NET_217, __A15_2__KY2RST, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15036(XT3_n, XB4_n, __A15_NET_220, GOJAM, DRPRST, __A15_1__DNRPTA, GND, DRPRST, XB0_n, XT4_n, __A15_1__KRPTA_n, __A15_NET_246, __A15_1__KRPTA_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15037(__A15_NET_294, __A15_NET_295, __A15_NET_242, __A15_NET_291, __A15_NET_241, __A15_NET_242, GND, __A15_NET_245, __A15_NET_237, __A15_NET_222, __A15_NET_213, __A15_NET_226, __A15_NET_216, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15038(__A15_NET_221, __A15_NET_214, __A15_NET_295, __A15_NET_239, __A15_NET_240, __A15_NET_242, GND, __A15_NET_290, __A15_NET_216, __A15_NET_214, __A15_1__PRPOR4, __A15_NET_296, __A15_1__PRPOR3, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U15039(__A15_NET_290, __A15_NET_232, __A15_NET_265, RL03_n, __A15_NET_297, RL04_n, GND, RL05_n, __A15_NET_298, RL02_n, __A15_NET_299, RL01_n, __A15_NET_310, p4VSW, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC27 U15040(__A15_NET_295, __A15_NET_243, __A15_NET_245, __A15_NET_234, __A15_NET_223, __A15_NET_221, GND, __A15_NET_224, __A15_NET_245, __A15_NET_225, __A15_NET_223, __A15_NET_244, __A15_NET_240, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U15041(__A15_NET_260, __A15_NET_221, __A15_NET_222, __A15_NET_216, __A15_NET_214,  , GND,  , __A15_2__RPTAD3, __A15_1__BBK3, CAD3, R6, __A15_NET_265, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15042(__A15_NET_213, __A15_NET_215, __A15_NET_213, __A15_NET_219, __A15_NET_217, __A15_NET_218, GND,  ,  ,  ,  , __A15_NET_214, __A15_NET_217, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15043(__A15_1__PRPOR2, __A15_1__PRPOR1, __A15_NET_220, __A15_2__RPTAD3, __A15_1__RRPA1_n, __A15_NET_229, GND, __A15_1__RRPA1_n, __A15_NET_232, __A15_2__RPTAD4, __A15_2__RPTAD4, CAD4, __A15_NET_297, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15044(RRPA, __A15_1__RRPA1_n, STRGAT, __A15_NET_227, __A15_1__F11, __A15_NET_228, GND, __A15_NET_272, __A15_1__F11_n, __A15_NET_273, S10, __A15_NET_271, S10_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15045(__A15_NET_298, __A15_2__RPTAD5, CAD5, __A15_2__RPTAD5, __A15_1__RRPA1_n, __A15_NET_260, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15046(CAD2, __A15_1__BBK2, CAD1, __A15_1__BBK1, RB1F, __A15_NET_310, GND, STR412, __A15_NET_227, __A15_NET_273, __A15_NET_228, __A15_NET_299, R6, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15047(__A15_NET_227, __A15_NET_271, __A15_NET_227, __A15_NET_273, __A15_NET_272, STR210, GND, STR19, __A15_NET_227, __A15_NET_271, __A15_NET_272, STR311, __A15_NET_228, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15048(__A15_NET_274, __A15_1__F16, __A15_1__F15, __A15_NET_269, __A15_1__F16, __A15_1__F15_n, GND, __A15_1__F15, __A15_1__F16_n, __A15_NET_287, __A15_2__NE036_n, __A15_1__F12, __A15_2__036L, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15049(__A15_NET_274, __A15_NET_268, __A15_1__F14_n, __A15_NET_270, __A15_1__F13_n, __A15_NET_285, GND, __A15_NET_282, __A15_1__F13, __A15_NET_284, __A15_1__F14, __A15_NET_283, __A15_NET_269, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15050(__A15_NET_268, __A15_NET_270, __A15_NET_268, __A15_NET_270, __A15_NET_282, __A15_2__NE01, GND, __A15_2__NE02, __A15_NET_268, __A15_NET_284, __A15_NET_285, __A15_2__NE00, __A15_NET_285, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15051(__A15_NET_268, __A15_NET_284, __A15_NET_283, __A15_NET_270, __A15_NET_285, __A15_2__NE04, GND, __A15_2__NE05, __A15_NET_283, __A15_NET_270, __A15_NET_282, __A15_2__NE03, __A15_NET_282, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15052(__A15_NET_283, __A15_NET_284, __A15_NET_283, __A15_NET_284, __A15_NET_282, __A15_2__NE07, GND, __A15_2__NE10, __A15_NET_286, __A15_NET_270, __A15_NET_285, __A15_2__NE06, __A15_NET_285, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15053(__A15_NET_287, __A15_NET_286, __A15_NET_251, STR14, __A15_2__NE012_n, ROPER, GND, LOMOD, __A15_NET_266, STR58, __A15_NET_267, ROPES, __A15_2__NE345_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15054(__A15_2__NE00, __A15_2__NE03, __A15_2__NE00, __A15_2__NE01, __A15_2__NE02, __A15_2__NE012_n, GND, __A15_2__NE147_n, __A15_2__NE01, __A15_2__NE04, __A15_2__NE07, __A15_2__NE036_n, __A15_2__NE06, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15055(__A15_2__NE04, __A15_2__NE03, __A15_2__NE02, __A15_2__NE05, __A15_2__NE10, __A15_2__NE2510_n, GND, __A15_2__NE6710_n, __A15_2__NE06, __A15_2__NE07, __A15_2__NE10, __A15_2__NE345_n, __A15_2__NE05, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15056(__A15_2__147H, __A15_2__NE147_n, __A15_1__F12_n, __A15_2__2510L, __A15_2__NE2510_n, __A15_1__F12, GND, __A15_2__NE036_n, __A15_1__F12_n, __A15_2__036H, __A15_2__NE147_n, __A15_1__F12, __A15_2__147L, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15057(__A15_2__2510H, __A15_2__NE2510_n, __A15_1__F12_n, __A15_NET_251, __A15_2__036L, __A15_2__147H, GND, __A15_2__2510L, __A15_2__036H, __A15_NET_267, __A15_2__147L, __A15_2__2510H, __A15_NET_262, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15058(__A15_2__036L, __A15_2__147L, __A15_2__147H, __A15_2__2510H, __A15_2__2510L, __A15_NET_261, GND,  ,  ,  ,  , __A15_NET_266, __A15_2__036H, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15059(__A15_NET_261, HIMOD, __A15_NET_262, STR912, __A15_2__NE6710_n, ROPET, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
endmodule