`include "components/agc_parts.v"

module timer(VCC, GND, SIM_RST, CLOCK, MSTRTP, MSTP, PHS2, PHS2_n, PHS3_n, PHS4, PHS4_n, RT, RT_n, WT, WT_n, CT, CT_n, CLK, TT_n, P01, P01_n, P02, P02_n, P03, P03_n, P04, P04_n, P05, P05_n, SBY, ALGA, STRT1, STRT2, GOJ1, STOPA, GOJAM, GOJAM_n, STOP, STOP_n, WL15, WL15_n, WL16, WL16_n, FS01_n, T01, T01_n, T02, T02_n, T03, T03_n, T04, T04_n, T05, T05_n, T06, T06_n, T07, T07_n, T08, T08_n, T09, T09_n, T10, T10_n, T11, T11_n, T12, T12_n, MONWT, Q2A, MGOJAM, MSTPIT_n);
    input wire SIM_RST;
    wire __A02_2__F01D;
    output wire PHS4;
    wire NET_175;
    wire NET_174;
    wire NET_173;
    wire __A02_2__F01A;
    wire __A02_2__F01B;
    output wire PHS2;
    wire __A02_3__OVF;
    wire __A02_3__UNF;
    wire NET_179;
    output wire P01_n;
    output wire WT;
    wire NET_172;
    output wire RT;
    output wire RT_n;
    output wire T03_n;
    wire NET_182;
    wire NET_180;
    output wire P05_n;
    wire NET_177;
    wire __A02_1__ovfstb_r4;
    output wire P03_n;
    wire __A02_1__ovfstb_r5;
    wire NET_164;
    wire __A02_1__RINGA_n;
    wire NET_166;
    wire NET_167;
    wire NET_160;
    wire NET_161;
    wire NET_162;
    wire NET_163;
    wire __A02_1__ODDSET_n;
    wire __A02_1__cdiv_2__FS_n;
    wire NET_168;
    wire NET_169;
    output wire T07;
    output wire T06;
    output wire T05;
    output wire T04;
    output wire T03;
    output wire T02;
    output wire T01;
    wire __A02_1__ovfstb_r2;
    wire __A02_1__ovfstb_r3;
    wire NET_171;
    wire __A02_1__ovfstb_r1;
    wire __A02_1__ovfstb_r6;
    output wire T09;
    output wire T08;
    wire __A02_3__T07DC_n;
    output wire T10_n;
    output wire P03;
    output wire P02;
    output wire P01;
    output wire T09_n;
    output wire P05;
    output wire P04;
    wire NET_170;
    input wire GOJ1;
    input wire WL16_n;
    wire NET_151;
    output wire Q2A;
    wire NET_153;
    wire NET_152;
    wire __A02_2__FS01;
    wire NET_154;
    wire NET_157;
    wire __A02_1__cdiv_1__B;
    wire NET_159;
    wire NET_158;
    output wire T10;
    output wire T11;
    output wire T12;
    wire __A02_3__T12DC_n;
    output wire P04_n;
    wire __A02_3__T04DC_n;
    wire __A02_3__T12SET;
    wire NET_149;
    output wire P02_n;
    wire __A02_1__RINGB_n;
    wire NET_147;
    wire NET_148;
    wire __A02_3__UNF_n;
    wire NET_146;
    wire NET_142;
    wire NET_144;
    wire NET_145;
    input wire MSTP;
    wire NET_143;
    wire NET_140;
    wire NET_141;
    wire __A02_3__OVF_n;
    wire __A02_3__MT09;
    wire NET_150;
    wire __A02_1__cdiv_1__D;
    wire NET_178;
    wire __A02_1__evnset;
    wire __A02_3__T02DC_n;
    input wire ALGA;
    output wire T11_n;
    wire __A02_3__MT05;
    wire __A02_3__T08DC_n;
    wire NET_139;
    wire NET_138;
    input wire CLOCK;
    wire NET_133;
    wire NET_132;
    wire NET_131;
    output wire STOP;
    wire NET_136;
    wire NET_135;
    wire NET_134;
    wire __A02_1__cdiv_2__D;
    wire __A02_1__cdiv_2__F;
    wire __A02_1__cdiv_2__A;
    wire __A02_1__cdiv_2__B;
    wire __A02_1__cdiv_2__C;
    wire __A02_1__cdiv_1__A;
    output wire T05_n;
    wire __A02_3__T06DC_n;
    wire __A02_3__T09DC_n;
    wire __A02_3__MT08;
    wire __A02_3__MT07;
    wire __A02_3__MT06;
    output wire PHS2_n;
    wire __A02_3__MT04;
    wire __A02_3__MT03;
    wire __A02_3__MT02;
    wire __A02_3__MT01;
    output wire GOJAM;
    wire __A02_1__cdiv_2__FS;
    wire NET_155;
    output wire CLK;
    output wire GOJAM_n;
    output wire T01_n;
    input wire WL15_n;
    wire NET_137;
    output wire PHS4_n;
    output wire T07_n;
    output wire STOPA;
    output wire FS01_n;
    output wire CT;
    wire __A02_3__MT10;
    wire __A02_3__MT11;
    wire __A02_3__MT12;
    input wire SBY;
    output wire CT_n;
    wire __A02_1__oddset;
    wire __A02_1__cdiv_1__FS_n;
    wire NET_165;
    output wire T12_n;
    input wire WL16;
    output wire MONWT;
    input wire WL15;
    input wire GND;
    wire NET_156;
    output wire T04_n;
    wire NET_117;
    input wire MSTRTP;
    wire __A02_1__cdiv_1__FS;
    input wire STRT1;
    input wire STRT2;
    output wire MGOJAM;
    wire __A02_3__T10DC_n;
    output wire T02_n;
    wire NET_181;
    input wire VCC;
    wire NET_176;
    output wire T08_n;
    output wire T06_n;
    output wire PHS3_n;
    output wire MSTPIT_n;
    wire __A02_1__EVNSET_n;
    wire __A02_3__T01DC_n;
    output wire TT_n;
    wire __A02_1__OVFSTB_n;
    output wire WT_n;
    wire __A02_2__F01C;
    wire __A02_3__T03DC_n;
    wire __A02_3__T05DC_n;
    output wire STOP_n;

    U74HC02 U9(__A02_1__ovfstb_r1, CT_n, __A02_1__ovfstb_r2, __A02_1__ovfstb_r2, __A02_1__ovfstb_r6, __A02_1__ovfstb_r1, GND, __A02_1__ovfstb_r4, __A02_1__ovfstb_r2, __A02_1__ovfstb_r3, __A02_1__ovfstb_r3, __A02_1__ovfstb_r1, __A02_1__ovfstb_r4, VCC, SIM_RST);
    U74HC04 U8(__A02_1__cdiv_2__D, __A02_1__RINGA_n, __A02_1__oddset, __A02_1__ODDSET_n, __A02_1__cdiv_2__C, __A02_1__RINGB_n, GND, __A02_1__evnset, __A02_1__RINGB_n, __A02_1__EVNSET_n, __A02_1__evnset, RT, __A02_1__cdiv_1__A, VCC, SIM_RST);
    U74HC04 U5(__A02_1__cdiv_1__FS_n, WT, WT, WT_n, WT, TT_n, GND, __A02_1__ovfstb_r5, __A02_1__ovfstb_r4, __A02_1__ovfstb_r6, __A02_1__ovfstb_r5, __A02_1__OVFSTB_n, __A02_1__ovfstb_r2, VCC, SIM_RST);
    wire U4_8_NC;
    wire U4_9_NC;
    wire U4_10_NC;
    wire U4_11_NC;
    wire U4_12_NC;
    wire U4_13_NC;
    U74HC02 U4(PHS4, __A02_1__cdiv_2__F, __A02_1__cdiv_1__A, __A02_1__oddset, STOP, __A02_1__RINGA_n, GND, U4_8_NC, U4_9_NC, U4_10_NC, U4_11_NC, U4_12_NC, U4_13_NC, VCC, SIM_RST);
    wire U7_8_NC;
    wire U7_9_NC;
    wire U7_10_NC;
    wire U7_11_NC;
    U74HC27 #(0, 1, 0) U7(__A02_1__cdiv_2__D, __A02_1__cdiv_2__F, __A02_1__cdiv_2__B, __A02_1__cdiv_2__F, __A02_1__cdiv_2__C, __A02_1__cdiv_2__A, GND, U7_8_NC, U7_9_NC, U7_10_NC, U7_11_NC, __A02_1__cdiv_2__B, __A02_1__cdiv_2__A, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U6(__A02_1__cdiv_2__D, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__FS, GND, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__A, __A02_1__cdiv_2__FS, __A02_1__cdiv_2__A, __A02_1__cdiv_2__FS, __A02_1__cdiv_2__C, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U1(__A02_1__cdiv_1__D, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__B, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__B, __A02_1__cdiv_1__FS, GND, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__A, __A02_1__cdiv_1__FS, __A02_1__cdiv_1__A, __A02_1__cdiv_1__FS, PHS2, VCC, SIM_RST);
    U74HC04 U3(__A02_1__cdiv_1__D, __A02_1__cdiv_2__F, PHS2, PHS2_n, PHS4, PHS4_n, GND, NET_117, __A02_1__cdiv_1__B, CT, NET_117, CT_n, CT, VCC, SIM_RST);
    wire U2_8_NC;
    wire U2_9_NC;
    wire U2_10_NC;
    wire U2_11_NC;
    U74HC27 #(0, 1, 0) U2(__A02_1__cdiv_1__D, CLOCK, __A02_1__cdiv_1__B, CLOCK, PHS2, __A02_1__cdiv_1__A, GND, U2_8_NC, U2_9_NC, U2_10_NC, U2_11_NC, __A02_1__cdiv_1__B, __A02_1__cdiv_1__A, VCC, SIM_RST);
    U74HC27 U19(SBY, ALGA, STRT1, STRT2, NET_134, NET_132, GND, NET_140, GND, NET_141, __A02_1__EVNSET_n, NET_131, MSTRTP, VCC, SIM_RST);
    wire U18_8_NC;
    wire U18_9_NC;
    wire U18_10_NC;
    wire U18_11_NC;
    U74HC27 #(0, 1, 0) U18(__A02_2__F01D, P01_n, __A02_2__F01B, P01_n, __A02_2__F01C, __A02_2__F01A, GND, U18_8_NC, U18_9_NC, U18_10_NC, U18_11_NC, __A02_2__F01B, __A02_2__F01A, VCC, SIM_RST);
    U74HC02 U35(T09, __A02_1__ODDSET_n, __A02_3__T09DC_n, NET_162, __A02_1__EVNSET_n, __A02_3__T09DC_n, GND, NET_181, NET_162, __A02_3__T10DC_n, __A02_1__EVNSET_n, NET_181, NET_160, VCC, SIM_RST);
    U74HC27 U34(GOJAM, NET_181, GOJAM, NET_178, __A02_3__T10DC_n, NET_181, GND, NET_178, GOJAM, NET_160, NET_163, NET_182, __A02_3__T09DC_n, VCC, SIM_RST);
    U74HC02 U33(__A02_3__T08DC_n, NET_179, NET_166, T08, __A02_1__EVNSET_n, __A02_3__T08DC_n, GND, __A02_1__ODDSET_n, __A02_3__T08DC_n, NET_159, NET_182, NET_159, __A02_3__T09DC_n, VCC, SIM_RST);
    U74HC02 U32(NET_167, __A02_1__ODDSET_n, __A02_3__T06DC_n, __A02_3__T07DC_n, NET_180, NET_167, GND, __A02_1__ODDSET_n, __A02_3__T07DC_n, T07, __A02_1__EVNSET_n, __A02_3__T07DC_n, NET_166, VCC, SIM_RST);
    U74HC27 U31(GOJAM, NET_180, GOJAM, NET_179, __A02_3__T07DC_n, NET_180, GND, NET_179, GOJAM, NET_182, __A02_3__T08DC_n, NET_173, __A02_3__T06DC_n, VCC, SIM_RST);
    U74HC02 U30(NET_155, __A02_3__T05DC_n, __A02_1__EVNSET_n, T05, __A02_3__T05DC_n, __A02_1__ODDSET_n, GND, NET_173, NET_155, __A02_3__T06DC_n, __A02_1__EVNSET_n, __A02_3__T06DC_n, T06, VCC, SIM_RST);
    U74HC27 U11(__A02_1__RINGB_n, P05_n, P04, P05, __A02_1__RINGA_n, NET_152, GND, NET_145, GND, NET_142, __A02_1__EVNSET_n, NET_151, P04_n, VCC, SIM_RST);
    wire U10_12_NC;
    wire U10_13_NC;
    U74HC04 U10(CT, PHS3_n, WT_n, CLK, WT_n, MONWT, GND, Q2A, WT_n, RT_n, RT, U10_12_NC, U10_13_NC, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U13(P02, NET_148, P02_n, P02_n, P02, NET_153, GND, __A02_1__RINGB_n, P02, NET_150, P02_n, __A02_1__RINGA_n, NET_149, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U12(P01, NET_151, P01_n, P01_n, P01, NET_152, GND, __A02_1__RINGA_n, P01, NET_148, P01_n, __A02_1__RINGB_n, NET_153, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U15(P04, NET_135, P04_n, P04_n, P04, NET_136, GND, __A02_1__RINGB_n, P04, NET_138, P04_n, __A02_1__RINGA_n, NET_137, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U14(P03, NET_150, P03_n, P03_n, P03, NET_149, GND, __A02_1__RINGA_n, P03, NET_135, P03_n, __A02_1__RINGB_n, NET_136, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U17(__A02_2__F01D, FS01_n, __A02_2__F01B, FS01_n, __A02_2__F01B, __A02_2__FS01, GND, FS01_n, __A02_2__F01A, __A02_2__FS01, __A02_2__F01A, __A02_2__FS01, __A02_2__F01C, VCC, SIM_RST);
    U74HC02 #(0, 1, 1, 0) U16(P05, NET_138, P05_n, P05_n, P05, NET_137, GND, NET_142, GOJ1, NET_134, __A02_1__EVNSET_n, NET_133, NET_146, VCC, SIM_RST);
    U74HC04 U43(T10, T10_n, T10_n, __A02_3__MT10, T11, T11_n, GND, __A02_3__MT11, T11_n, T12_n, T12, __A02_3__MT12, T12_n, VCC, SIM_RST);
    wire U39_10_NC;
    wire U39_11_NC;
    wire U39_12_NC;
    wire U39_13_NC;
    U74LVC07 U39(NET_154, __A02_3__T12SET, NET_156, __A02_3__T12SET, NET_158, __A02_3__T12SET, GND, __A02_3__T12SET, NET_157, U39_10_NC, U39_11_NC, U39_12_NC, U39_13_NC, VCC, SIM_RST);
    U74HC27 U38(NET_172, NET_171, NET_182, NET_181, __A02_1__EVNSET_n, NET_158, GND, NET_157, NET_173, NET_180, NET_179, NET_156, NET_175, VCC, SIM_RST);
    wire U44_8_NC;
    wire U44_9_NC;
    wire U44_10_NC;
    wire U44_11_NC;
    U74HC27 U44(WL15_n, WL16, __A02_1__OVFSTB_n, WL15, WL16_n, __A02_3__UNF, GND, U44_8_NC, U44_9_NC, U44_10_NC, U44_11_NC, __A02_3__OVF, __A02_1__OVFSTB_n, VCC, SIM_RST);
    pullup R1(NET_142);
    pullup R2(__A02_3__T12SET);
    U74HC27 U24(__A02_3__T12SET, GOJAM, __A02_3__T01DC_n, NET_177, GOJAM, NET_174, GND, NET_177, __A02_3__T02DC_n, NET_175, GOJAM, __A02_3__T12DC_n, NET_176, VCC, SIM_RST);
    U74HC02 U25(NET_176, __A02_3__T12DC_n, NET_174, NET_164, __A02_3__T12DC_n, __A02_1__ODDSET_n, GND, __A02_3__T12DC_n, __A02_1__EVNSET_n, T12, NET_164, NET_174, __A02_3__T01DC_n, VCC, SIM_RST);
    U74HC02 U26(NET_169, __A02_3__T01DC_n, __A02_1__EVNSET_n, T01, __A02_3__T01DC_n, __A02_1__ODDSET_n, GND, NET_169, NET_177, __A02_3__T02DC_n, __A02_3__T02DC_n, __A02_1__ODDSET_n, NET_168, VCC, SIM_RST);
    U74HC02 U27(T02, __A02_3__T02DC_n, __A02_1__EVNSET_n, __A02_3__T03DC_n, NET_168, NET_175, GND, __A02_3__T03DC_n, __A02_1__EVNSET_n, NET_170, __A02_3__T03DC_n, __A02_1__ODDSET_n, T03, VCC, SIM_RST);
    wire U20_5_NC;
    wire U20_6_NC;
    wire U20_8_NC;
    wire U20_9_NC;
    wire U20_10_NC;
    wire U20_11_NC;
    wire U20_12_NC;
    wire U20_13_NC;
    U74LVC07 U20(NET_131, NET_142, NET_132, NET_142, U20_5_NC, U20_6_NC, GND, U20_8_NC, U20_9_NC, U20_10_NC, U20_11_NC, U20_12_NC, U20_13_NC, VCC, SIM_RST);
    U74HC04 U21(NET_142, NET_133, MSTP, NET_141, GOJAM_n, GOJAM, GND, MGOJAM, GOJAM, STOP, STOP_n, MSTPIT_n, STOP, VCC, SIM_RST);
    wire U22_11_NC;
    wire U22_12_NC;
    wire U22_13_NC;
    U74HC02 U22(NET_139, __A02_1__EVNSET_n, MSTP, GOJAM_n, STRT2, STOPA, GND, STOPA, NET_143, STOP_n, U22_11_NC, U22_12_NC, U22_13_NC, VCC, SIM_RST);
    U74HC02 #(1, 0, 1, 0) U23(NET_144, NET_145, STOPA, STOPA, NET_144, NET_146, GND, NET_140, NET_143, NET_147, NET_147, NET_139, NET_143, VCC, SIM_RST);
    wire U45_5_NC;
    wire U45_6_NC;
    wire U45_8_NC;
    wire U45_9_NC;
    wire U45_10_NC;
    wire U45_11_NC;
    wire U45_12_NC;
    wire U45_13_NC;
    U74HC04 U45(__A02_3__OVF, __A02_3__OVF_n, __A02_3__UNF, __A02_3__UNF_n, U45_5_NC, U45_6_NC, GND, U45_8_NC, U45_9_NC, U45_10_NC, U45_11_NC, U45_12_NC, U45_13_NC, VCC, SIM_RST);
    U74HC27 U28(__A02_3__T03DC_n, NET_171, __A02_3__T04DC_n, NET_172, GOJAM, NET_171, GND, NET_172, __A02_3__T05DC_n, NET_173, GOJAM, NET_175, GOJAM, VCC, SIM_RST);
    U74HC02 U29(__A02_3__T04DC_n, NET_170, NET_171, NET_165, __A02_3__T04DC_n, __A02_1__ODDSET_n, GND, __A02_3__T04DC_n, __A02_1__EVNSET_n, T04, NET_165, NET_172, __A02_3__T05DC_n, VCC, SIM_RST);
    wire U37_4_NC;
    wire U37_5_NC;
    wire U37_6_NC;
    wire U37_8_NC;
    wire U37_9_NC;
    wire U37_10_NC;
    wire U37_11_NC;
    wire U37_12_NC;
    wire U37_13_NC;
    U74HC02 U37(NET_154, NET_177, NET_174, U37_4_NC, U37_5_NC, U37_6_NC, GND, U37_8_NC, U37_9_NC, U37_10_NC, U37_11_NC, U37_12_NC, U37_13_NC, VCC, SIM_RST);
    U74HC02 U36(NET_161, __A02_1__ODDSET_n, __A02_3__T10DC_n, NET_163, NET_178, NET_161, GND, __A02_1__EVNSET_n, __A02_3__T10DC_n, T10, __A02_1__ODDSET_n, NET_163, T11, VCC, SIM_RST);
    U74HC04 U40(T01, T01_n, T01_n, __A02_3__MT01, T02, T02_n, GND, __A02_3__MT02, T02_n, T03_n, T03, __A02_3__MT03, T03_n, VCC, SIM_RST);
    U74HC04 U41(T04, T04_n, T04_n, __A02_3__MT04, T05, T05_n, GND, __A02_3__MT05, T05_n, T06_n, T06, __A02_3__MT06, T06_n, VCC, SIM_RST);
    U74HC04 U42(T07, T07_n, T07_n, __A02_3__MT07, T08, T08_n, GND, __A02_3__MT08, T08_n, T09_n, T09, __A02_3__MT09, T09_n, VCC, SIM_RST);
endmodule