`timescale 1ns/1ps

module fpga_agc(VCC, GND, SIM_RST, SIM_CLK, ALGA, C24A, C25A, C26A, C27A, C30A, C37P, C40P, C41P, C42P, C43P, C44P, CDUSTB_n, CH01, CH02, CH03, CH04, CH05, CH06, CH07, CH08, CH09, CH10, CH11, CH12, CH13, CH14, CH16, CHINC_n, CLOCK, DINC, DINC_n, FETCH0, FETCH0_n, FETCH1, G16SW_n, INCSET_n, INKL, INKL_n, INOTLD, MCDU, MDT01, MDT02, MDT03, MDT04, MDT05, MDT06, MDT07, MDT08, MDT09, MDT10, MDT11, MDT12, MDT13, MDT14, MDT15, MDT16, MINC, MNHRPT, MONPAR, MONPCH, MONWBK, MON_n, MSTP, MSTRTP, MTCSAI, OVNHRP, PCDU, PIPPLS_n, RCHAT_n, RCHBT_n, RUPTOR_n, SA01, SA02, SA03, SA04, SA05, SA06, SA07, SA08, SA09, SA10, SA11, SA12, SA13, SA14, SA16, SAP, SBY, SHANC_n, SHIFT, SHIFT_n, STBE, STBF, STFET1_n, STORE1_n, STRT1, STRT2, TPARG_n, XB0_n, XB1_n, XB2_n, XB3_n, XB4_n, XB5_n, XB6_n, XB7_n, XT0_n, XT1_n, XT2_n, XT3_n, XT4_n, XT5_n, XT6_n, YB0_n, YT0_n, MGOJAM, MT01, MT02, MT03, MT04, MT05, MT06, MT07, MT08, MT09, MT10, MT11, MT12);

    input wire VCC;
    input wire GND;
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire ALGA;
    input wire C24A;
    input wire C25A;
    input wire C26A;
    input wire C27A;
    input wire C30A;
    input wire C37P;
    input wire C40P;
    input wire C41P;
    input wire C42P;
    input wire C43P;
    input wire C44P;
    input wire CDUSTB_n;
    input wire CH01;
    input wire CH02;
    input wire CH03;
    input wire CH04;
    input wire CH05;
    input wire CH06;
    input wire CH07;
    input wire CH08;
    input wire CH09;
    input wire CH10;
    input wire CH11;
    input wire CH12;
    input wire CH13;
    input wire CH14;
    input wire CH16;
    input wire CHINC_n;
    input wire CLOCK;
    input wire DINC;
    input wire DINC_n;
    input wire FETCH0;
    input wire FETCH0_n;
    input wire FETCH1;
    input wire G16SW_n;
    input wire INCSET_n;
    input wire INKL;
    input wire INKL_n;
    input wire INOTLD;
    input wire MCDU;
    input wire MDT01;
    input wire MDT02;
    input wire MDT03;
    input wire MDT04;
    input wire MDT05;
    input wire MDT06;
    input wire MDT07;
    input wire MDT08;
    input wire MDT09;
    input wire MDT10;
    input wire MDT11;
    input wire MDT12;
    input wire MDT13;
    input wire MDT14;
    input wire MDT15;
    input wire MDT16;
    input wire MINC;
    input wire MNHRPT;
    input wire MONPAR;
    input wire MONPCH;
    input wire MONWBK;
    input wire MON_n;
    input wire MSTP;
    input wire MSTRTP;
    input wire MTCSAI;
    input wire OVNHRP;
    input wire PCDU;
    input wire PIPPLS_n;
    input wire RCHAT_n;
    input wire RCHBT_n;
    input wire RUPTOR_n;
    input wire SA01;
    input wire SA02;
    input wire SA03;
    input wire SA04;
    input wire SA05;
    input wire SA06;
    input wire SA07;
    input wire SA08;
    input wire SA09;
    input wire SA10;
    input wire SA11;
    input wire SA12;
    input wire SA13;
    input wire SA14;
    input wire SA16;
    input wire SAP;
    input wire SBY;
    input wire SHANC_n;
    input wire SHIFT;
    input wire SHIFT_n;
    input wire STBE;
    input wire STBF;
    input wire STFET1_n;
    input wire STORE1_n;
    input wire STRT1;
    input wire STRT2;
    input wire TPARG_n;
    input wire XB0_n;
    input wire XB1_n;
    input wire XB2_n;
    input wire XB3_n;
    input wire XB4_n;
    input wire XB5_n;
    input wire XB6_n;
    input wire XB7_n;
    input wire XT0_n;
    input wire XT1_n;
    input wire XT2_n;
    input wire XT3_n;
    input wire XT4_n;
    input wire XT5_n;
    input wire XT6_n;
    input wire YB0_n;
    input wire YT0_n;
    output wire MGOJAM;
    output wire MT01;
    output wire MT02;
    output wire MT03;
    output wire MT04;
    output wire MT05;
    output wire MT06;
    output wire MT07;
    output wire MT08;
    output wire MT09;
    output wire MT10;
    output wire MT11;
    output wire MT12;
    wire A2XG_n;
    wand A2X_n;
    wire A2X_n_U5012_10;
    wire A2X_n_U5046_8;
    wire A2X_n_U6004_6;
    wire AD0;
    wire ADS0;
    wire AUG0_n;
    wire B15X;
    wire BR1;
    wire BR12B_n;
    wire BR1B2B;
    wire BR1B2B_n;
    wire BR1B2_n;
    wire BR1_n;
    wire BR2;
    wire BR2_n;
    wire BRDIF_n;
    wire BXVX;
    wire CAG;
    wire CBG;
    wire CCS0;
    wire CCS0_n;
    wire CGG;
    wire CGMC;
    wire CI01_n;
    wire CI05_n;
    wire CI09_n;
    wire CI13_n;
    wand CI_n;
    wire CI_n_U4061_12;
    wire CI_n_U5018_2;
    wire CI_n_U5046_10;
    wire CI_n_U6047_2;
    wire CLG1G;
    wire CLG2G;
    wire CLK;
    wire CLXC;
    wand CO06;
    wire CO06_U8041_2;
    wire CO06_U8050_2;
    wand CO10;
    wire CO10_U9041_2;
    wire CO10_U9050_2;
    wand CO14;
    wire CO14_U10041_2;
    wire CO14_U10050_2;
    wire CQG;
    wire CSG;
    wire CT;
    wire CT_n;
    wire CUG;
    wire CYL_n;
    wire CYR_n;
    wire CZG;
    wire DAS0;
    wire DAS0_n;
    wire DAS1;
    wire DAS1_n;
    wire DCA0;
    wire DCS0;
    wire DIM0_n;
    wire DIVSTG;
    wire DIV_n;
    wire DV1;
    wire DV1376;
    wire DV1376_n;
    wire DV1_n;
    wire DV376_n;
    wire DV4;
    wire DV4B1B;
    wire DV4_n;
    wire DVST;
    wire DXCH0;
    wire EAC_n;
    wire EDOP_n;
    wire EXST0_n;
    wire EXST1_n;
    wire EXT;
    wire EXTPLS;
    wire FS01_n;
    wire FUTEXT;
    wire G01;
    wire G01ED;
    wand G01_n;
    wire G01_n_U8013_6;
    wire G01_n_U8013_8;
    wire G02;
    wire G02ED;
    wire G03;
    wire G03ED;
    wire G04;
    wire G04ED;
    wire G05;
    wire G05ED;
    wand G05_n;
    wire G05_n_U9013_6;
    wire G05_n_U9013_8;
    wire G06;
    wire G06ED;
    wand G06_n;
    wire G06_n_U9028_10;
    wire G06_n_U9028_12;
    wire G07;
    wire G07ED;
    wand G07_n;
    wire G07_n_U9050_6;
    wire G07_n_U9050_8;
    wire G08;
    wire G09;
    wand G09_n;
    wire G09_n_U10013_6;
    wire G09_n_U10013_8;
    wire G10;
    wand G10_n;
    wire G10_n_U10028_10;
    wire G10_n_U10028_12;
    wire G11;
    wand G11_n;
    wire G11_n_U10050_6;
    wire G11_n_U10050_8;
    wire G12;
    wire G13;
    wand G13_n;
    wire G13_n_U11013_6;
    wire G13_n_U11013_8;
    wire G14;
    wand G14_n;
    wire G14_n_U11028_10;
    wire G14_n_U11028_12;
    wire G15;
    wand G15_n;
    wire G15_n_U11050_6;
    wire G15_n_U11050_8;
    wire G16;
    wire G2LSG_n;
    wire GEQZRO_n;
    wire GINH;
    wire GOJ1;
    wire GOJ1_n;
    wire GOJAM;
    wire GOJAM_n;
    wire IC1;
    wire IC10;
    wire IC10_n;
    wire IC11;
    wire IC11_n;
    wire IC12;
    wire IC12_n;
    wire IC13;
    wire IC14;
    wire IC15;
    wire IC15_n;
    wire IC16;
    wire IC16_n;
    wire IC17;
    wire IC2;
    wire IC2_n;
    wire IC3;
    wire IC4;
    wire IC5;
    wire IC5_n;
    wire IC6;
    wire IC7;
    wire IC8_n;
    wire IC9;
    wire INCR0;
    wand INHPLS;
    wire INHPLS_U12016_10;
    wire INHPLS_U12016_12;
    wire INOUT;
    wire INOUT_n;
    wire KRPT;
    wand L01_n;
    wire L01_n_U8007_6;
    wand L02_n;
    wire L02_n_U8013_12;
    wand L04_n;
    wire L04_n_U8050_12;
    wand L08_n;
    wire L08_n_U9050_12;
    wand L12_n;
    wire L12_n_U10050_12;
    wand L15_n;
    wire L15_n_U11041_6;
    wire L2GDG_n;
    wire L2GD_n;
    wire MASK0;
    wire MASK0_n;
    wire MCRO_n;
    wire MONEX;
    wand MONEX_n;
    wire MONEX_n_U5005_2;
    wire MONEX_n_U6029_6;
    wire MONWT;
    wire MP0;
    wire MP0T10;
    wire MP0_n;
    wire MP1;
    wire MP1_n;
    wire MP3;
    wire MP3A;
    wire MP3_n;
    wire MSTPIT_n;
    wire MSU0;
    wire MSU0_n;
    wire NDR100_n;
    wire NDX0_n;
    wire NDXX1_n;
    wire NEAC;
    wire NISQ;
    wire OCTAD2;
    wire OVF_n;
    wire P01;
    wire P01_n;
    wire P02;
    wire P02_n;
    wire P03;
    wire P03_n;
    wire P04;
    wire P04_n;
    wire P05;
    wire P05_n;
    wire PHS2;
    wire PHS2_n;
    wire PHS3_n;
    wire PHS4;
    wire PHS4_n;
    wire PIFL_n;
    wire PINC;
    wire PONEX;
    wire PRINC;
    wire PTWOX;
    wire Q2A;
    wire QC0_n;
    wire QC1_n;
    wire QC2_n;
    wire QC3_n;
    wire QXCH0_n;
    wire R15;
    wire R1C;
    wand R1C_n;
    wire R1C_n_U4063_10;
    wire R1C_n_U6029_12;
    wire R6;
    wire RAD;
    wire RADRG;
    wire RADRZ;
    wire RAG_n;
    wire RAND0;
    wand RA_n;
    wire RA_n_U4039_10;
    wire RA_n_U4045_8;
    wire RA_n_U5005_8;
    wire RA_n_U5024_4;
    wire RA_n_U5041_12;
    wire RB1;
    wand RB1_n;
    wire RB1_n_U4063_6;
    wire RB1_n_U6029_10;
    wire RB2;
    wire RBHG_n;
    wire RBLG_n;
    wire RBSQ;
    wand RB_n;
    wire RB_n_U4039_2;
    wire RB_n_U4061_10;
    wire RB_n_U5005_6;
    wire RB_n_U5018_10;
    wire RB_n_U5051_2;
    wire RB_n_U6004_8;
    wire RB_n_U6037_8;
    wire RCG_n;
    wire RCH_n;
    wand RC_n;
    wire RC_n_U4039_4;
    wire RC_n_U4061_8;
    wire RC_n_U5012_8;
    wire RC_n_U5024_10;
    wire RC_n_U5051_10;
    wire RC_n_U6047_6;
    wire RC_n_U6052_8;
    wire READ0;
    wand RELPLS;
    wire RELPLS_U12016_6;
    wire RELPLS_U12016_8;
    wire RGG_n;
    wand RG_n;
    wire RG_n_U5012_6;
    wire RG_n_U5046_2;
    wire RG_n_U5046_4;
    wire RG_n_U5061_10;
    wire RG_n_U6014_8;
    wire RL10BB;
    wire RLG_n;
    wand RL_n;
    wire RL_n_U5005_12;
    wire RL_n_U5041_10;
    wire ROR0;
    wand RPTSET;
    wire RPTSET_U3011_2;
    wire RPTSET_U3011_4;
    wire RPTSET_U3011_6;
    wire RPTSET_U6052_4;
    wire RQG_n;
    wire RQ_n;
    wire RRPA;
    wire RSC_n;
    wire RSM3;
    wire RSM3_n;
    wire RSTSTG;
    wire RT;
    wire RT_n;
    wire RUG_n;
    wire RULOG_n;
    wire RUPT0;
    wire RUPT1;
    wire RUS_n;
    wand RU_n;
    wire RU_n_U5024_2;
    wire RU_n_U5061_4;
    wire RU_n_U5061_6;
    wire RU_n_U6014_12;
    wire RU_n_U6037_2;
    wire RU_n_U6052_6;
    wire RXOR0;
    wire RXOR0_n;
    wire RZG_n;
    wand RZ_n;
    wire RZ_n_U5005_4;
    wire RZ_n_U5018_4;
    wire RZ_n_U5051_4;
    wire RZ_n_U6052_2;
    wire S11;
    wire S12;
    wire SB2_n;
    wand SCAD;
    wire SCAD_U5051_6;
    wire SCAD_U5051_8;
    wire SCAD_n;
    wire SQ0_n;
    wire SQ1_n;
    wire SQ2_n;
    wire SQEXT_n;
    wire SQR10;
    wire SQR10_n;
    wire SQR12_n;
    wire SR_n;
    wire ST0_n;
    wire ST1;
    wire ST1_n;
    wire ST2;
    wand ST2_n;
    wire ST2_n_U5024_6;
    wire ST2_n_U6047_12;
    wire ST3_n;
    wire STD2;
    wire STOP;
    wire STOPA;
    wire STOP_n;
    wire STRTFC;
    wire SU0;
    wire SUMA15_n;
    wire SUMA16_n;
    wire SUMB15_n;
    wire SUMB16_n;
    wire T01;
    wire T01_n;
    wire T02;
    wire T02_n;
    wire T03;
    wire T03_n;
    wire T04;
    wire T04_n;
    wire T05;
    wire T05_n;
    wire T06;
    wire T06_n;
    wire T07;
    wire T07_n;
    wire T08;
    wire T08_n;
    wire T09;
    wire T09_n;
    wire T10;
    wire T10_n;
    wire T11;
    wire T11_n;
    wire T12;
    wire T12A;
    wire T12USE_n;
    wire T12_n;
    wire TC0;
    wire TC0_n;
    wire TCF0;
    wire TCSAJ3_n;
    wire TL15;
    wand TMZ_n;
    wire TMZ_n_U4045_12;
    wire TMZ_n_U5012_2;
    wire TMZ_n_U5067_6;
    wand TOV_n;
    wire TOV_n_U5061_2;
    wire TOV_n_U6019_4;
    wire TPZG_n;
    wire TRSM;
    wire TS0;
    wire TS0_n;
    wand TSGN_n;
    wire TSGN_n_U4063_2;
    wire TSGN_n_U4063_4;
    wire TSGN_n_U5061_12;
    wire TSGN_n_U5067_10;
    wire TSGU_n;
    wire TSUDO_n;
    wire TT_n;
    wire TWOX;
    wire U2BBK;
    wire UNF_n;
    wire US2SG;
    wire WAG_n;
    wire WALSG_n;
    wire WAND0;
    wand WA_n;
    wire WA_n_U5005_10;
    wire WA_n_U5024_12;
    wire WA_n_U5058_6;
    wire WA_n_U6029_8;
    wire WA_n_U6047_4;
    wire WBG_n;
    wand WB_n;
    wire WB_n_U5018_12;
    wire WB_n_U5041_2;
    wire WB_n_U5041_4;
    wire WB_n_U5061_8;
    wire WB_n_U6014_10;
    wire WCH_n;
    wire WEDOPG_n;
    wire WG1G_n;
    wire WG2G_n;
    wire WG3G_n;
    wire WG4G_n;
    wire WG5G_n;
    wand WG_n;
    wire WG_n_U4039_12;
    wire WG_n_U4045_10;
    wire WG_n_U4045_2;
    wire WG_n_U5012_4;
    wire WG_n_U6019_8;
    wire WG_n_U6037_6;
    wire WHOMP;
    wire WHOMPA;
    wire WL01_n;
    wire WL02_n;
    wire WL03_n;
    wire WL04_n;
    wire WL05_n;
    wire WL06_n;
    wire WL07_n;
    wire WL08_n;
    wire WL09_n;
    wire WL10_n;
    wire WL11_n;
    wire WL12_n;
    wire WL13_n;
    wire WL14_n;
    wire WL15;
    wire WL15_n;
    wire WL16;
    wire WL16_n;
    wire WLG_n;
    wand WL_n;
    wire WL_n_U4061_6;
    wire WL_n_U5067_4;
    wire WL_n_U6014_6;
    wire WOR0;
    wire WQG_n;
    wire WQ_n;
    wand WSC_n;
    wire WSC_n_U6019_6;
    wire WSC_n_U6037_4;
    wire WSG_n;
    wand WS_n;
    wire WS_n_U5035_12;
    wire WS_n_U6041_8;
    wire WT;
    wire WT_n;
    wand WY12_n;
    wire WY12_n_U5018_6;
    wire WY12_n_U5046_12;
    wire WYDG_n;
    wire WYDLOG_n;
    wand WYD_n;
    wire WYD_n_U5067_8;
    wire WYD_n_U6004_10;
    wire WYHIG_n;
    wire WYLOG_n;
    wand WY_n;
    wire WY_n_U4061_2;
    wire WY_n_U4061_4;
    wire WY_n_U5012_12;
    wire WY_n_U5024_8;
    wire WY_n_U5046_6;
    wire WY_n_U6004_12;
    wire WZG_n;
    wand WZ_n;
    wire WZ_n_U5018_8;
    wire WZ_n_U5058_12;
    wire WZ_n_U6019_2;
    wire XUY01_n;
    wire XUY02_n;
    wire XUY05_n;
    wire XUY06_n;
    wire XUY09_n;
    wire XUY10_n;
    wire XUY13_n;
    wire XUY14_n;
    wire ZAP_n;
    wire __A01_1__CHAT01;
    wire __A01_1__CHAT02;
    wire __A01_1__CHAT03;
    wire __A01_1__CHAT04;
    wire __A01_1__CHAT05;
    wire __A01_1__CHAT06;
    wire __A01_1__CHAT07;
    wire __A01_1__CHAT08;
    wire __A01_1__CHAT09;
    wire __A01_1__CHAT10;
    wire __A01_1__CHAT11;
    wire __A01_1__CHAT12;
    wire __A01_1__F02A;
    wire __A01_1__F02B;
    wire __A01_1__F03A;
    wire __A01_1__F03B;
    wire __A01_1__F04A;
    wire __A01_1__F04B;
    wire __A01_1__F05A;
    wire __A01_1__F05B;
    wire __A01_1__F06A;
    wire __A01_1__F06B;
    wire __A01_1__F07A;
    wire __A01_1__F07B;
    wire __A01_1__F08A;
    wire __A01_1__F08B;
    wire __A01_1__F09A;
    wire __A01_1__F09B;
    wire __A01_1__F10A;
    wire __A01_1__F10B;
    wire __A01_1__F11A;
    wire __A01_1__F11B;
    wire __A01_1__F12A;
    wire __A01_1__F12B;
    wire __A01_1__F13A;
    wire __A01_1__F13B;
    wire __A01_1__F14A;
    wire __A01_1__F14B;
    wire __A01_1__F15A;
    wire __A01_1__F15B;
    wire __A01_1__F16A;
    wire __A01_1__F16B;
    wire __A01_1__F17A;
    wire __A01_1__F17B;
    wire __A01_1__FS02;
    wire __A01_1__FS02A;
    wire __A01_1__FS03;
    wire __A01_1__FS03A;
    wire __A01_1__FS04;
    wire __A01_1__FS04A;
    wire __A01_1__FS05;
    wire __A01_1__FS05A;
    wire __A01_1__FS06;
    wire __A01_1__FS07;
    wire __A01_1__FS08;
    wire __A01_1__FS09;
    wire __A01_1__FS10;
    wire __A01_1__FS11;
    wire __A01_1__FS12;
    wire __A01_1__FS13;
    wire __A01_1__FS14;
    wire __A01_1__FS15;
    wire __A01_1__FS16;
    wire __A01_1__FS17;
    wire __A01_1__scaler_s10__FS_n;
    wire __A01_1__scaler_s11__FS_n;
    wire __A01_1__scaler_s12__FS_n;
    wire __A01_1__scaler_s13__FS_n;
    wire __A01_1__scaler_s14__FS_n;
    wire __A01_1__scaler_s15__FS_n;
    wire __A01_1__scaler_s16__FS_n;
    wire __A01_1__scaler_s17__FS_n;
    wire __A01_1__scaler_s2__FS_n;
    wire __A01_1__scaler_s3__FS_n;
    wire __A01_1__scaler_s4__FS_n;
    wire __A01_1__scaler_s5__FS_n;
    wire __A01_1__scaler_s6__FS_n;
    wire __A01_1__scaler_s7__FS_n;
    wire __A01_1__scaler_s8__FS_n;
    wire __A01_1__scaler_s9__FS_n;
    wire __A01_2__CHAT13;
    wire __A01_2__CHAT14;
    wire __A01_2__CHBT01;
    wire __A01_2__CHBT02;
    wire __A01_2__CHBT03;
    wire __A01_2__CHBT04;
    wire __A01_2__CHBT05;
    wire __A01_2__CHBT06;
    wire __A01_2__CHBT07;
    wire __A01_2__CHBT08;
    wire __A01_2__CHBT09;
    wire __A01_2__CHBT10;
    wire __A01_2__CHBT11;
    wire __A01_2__CHBT12;
    wire __A01_2__CHBT13;
    wire __A01_2__CHBT14;
    wire __A01_2__F18A;
    wire __A01_2__F18B;
    wire __A01_2__F19A;
    wire __A01_2__F19B;
    wire __A01_2__F20A;
    wire __A01_2__F20B;
    wire __A01_2__F21A;
    wire __A01_2__F21B;
    wire __A01_2__F22A;
    wire __A01_2__F22B;
    wire __A01_2__F23A;
    wire __A01_2__F23B;
    wire __A01_2__F24A;
    wire __A01_2__F24B;
    wire __A01_2__F25A;
    wire __A01_2__F25B;
    wire __A01_2__F26A;
    wire __A01_2__F26B;
    wire __A01_2__F27A;
    wire __A01_2__F27B;
    wire __A01_2__F28A;
    wire __A01_2__F28B;
    wire __A01_2__F29A;
    wire __A01_2__F29B;
    wire __A01_2__F30A;
    wire __A01_2__F30B;
    wire __A01_2__F31A;
    wire __A01_2__F31B;
    wire __A01_2__F32A;
    wire __A01_2__F32B;
    wire __A01_2__F33A;
    wire __A01_2__F33B;
    wire __A01_2__FS18;
    wire __A01_2__FS19;
    wire __A01_2__FS20;
    wire __A01_2__FS21;
    wire __A01_2__FS22;
    wire __A01_2__FS23;
    wire __A01_2__FS24;
    wire __A01_2__FS25;
    wire __A01_2__FS26;
    wire __A01_2__FS27;
    wire __A01_2__FS28;
    wire __A01_2__FS29;
    wire __A01_2__FS30;
    wire __A01_2__FS31;
    wire __A01_2__FS32;
    wire __A01_2__FS33;
    wire __A01_2__scaler_s18__FS_n;
    wire __A01_2__scaler_s19__FS_n;
    wire __A01_2__scaler_s20__FS_n;
    wire __A01_2__scaler_s21__FS_n;
    wire __A01_2__scaler_s22__FS_n;
    wire __A01_2__scaler_s23__FS_n;
    wire __A01_2__scaler_s24__FS_n;
    wire __A01_2__scaler_s25__FS_n;
    wire __A01_2__scaler_s26__FS_n;
    wire __A01_2__scaler_s27__FS_n;
    wire __A01_2__scaler_s28__FS_n;
    wire __A01_2__scaler_s29__FS_n;
    wire __A01_2__scaler_s30__FS_n;
    wire __A01_2__scaler_s31__FS_n;
    wire __A01_2__scaler_s32__FS_n;
    wire __A01_2__scaler_s33__FS_n;
    wire __A01_NET_143;
    wire __A01_NET_155;
    wire __A01_NET_168;
    wire __A01_NET_169;
    wire __A01_NET_170;
    wire __A01_NET_171;
    wire __A01_NET_172;
    wire __A01_NET_173;
    wire __A01_NET_174;
    wire __A01_NET_175;
    wire __A01_NET_176;
    wire __A01_NET_177;
    wire __A01_NET_178;
    wire __A01_NET_179;
    wire __A01_NET_180;
    wire __A01_NET_181;
    wire __A01_NET_182;
    wire __A01_NET_183;
    wire __A01_NET_184;
    wire __A01_NET_185;
    wire __A01_NET_186;
    wire __A01_NET_187;
    wire __A01_NET_188;
    wire __A01_NET_189;
    wire __A01_NET_190;
    wire __A01_NET_191;
    wire __A01_NET_192;
    wire __A01_NET_193;
    wire __A01_NET_194;
    wire __A01_NET_195;
    wire __A01_NET_196;
    wire __A01_NET_197;
    wire __A01_NET_198;
    wire __A01_NET_199;
    wire __A01_NET_200;
    wire __A01_NET_201;
    wire __A01_NET_202;
    wire __A01_NET_203;
    wire __A01_NET_204;
    wire __A01_NET_205;
    wire __A01_NET_206;
    wire __A01_NET_207;
    wire __A01_NET_208;
    wire __A01_NET_209;
    wire __A01_NET_210;
    wire __A01_NET_211;
    wire __A01_NET_212;
    wire __A01_NET_213;
    wire __A01_NET_214;
    wire __A01_NET_215;
    wire __A01_NET_216;
    wire __A01_NET_217;
    wire __A01_NET_218;
    wire __A01_NET_219;
    wire __A01_NET_220;
    wire __A01_NET_221;
    wire __A01_NET_222;
    wire __A01_NET_223;
    wire __A01_NET_224;
    wire __A01_NET_225;
    wire __A01_NET_226;
    wire __A01_NET_227;
    wire __A01_NET_228;
    wire __A01_NET_229;
    wire __A01_NET_230;
    wire __A01_NET_231;
    wire __A02_1__EVNSET_n;
    wire __A02_1__ODDSET_n;
    wire __A02_1__OVFSTB_n;
    wire __A02_1__RINGA_n;
    wire __A02_1__RINGB_n;
    wire __A02_1__cdiv_1__A;
    wire __A02_1__cdiv_1__B;
    wire __A02_1__cdiv_1__D;
    wire __A02_1__cdiv_1__FS;
    wire __A02_1__cdiv_1__FS_n;
    wire __A02_1__cdiv_2__A;
    wire __A02_1__cdiv_2__B;
    wire __A02_1__cdiv_2__C;
    wire __A02_1__cdiv_2__D;
    wire __A02_1__cdiv_2__F;
    wire __A02_1__cdiv_2__FS;
    wire __A02_1__cdiv_2__FS_n;
    wire __A02_1__evnset;
    wire __A02_1__oddset;
    wire __A02_1__ovfstb_r1;
    wire __A02_1__ovfstb_r2;
    wire __A02_1__ovfstb_r3;
    wire __A02_1__ovfstb_r4;
    wire __A02_1__ovfstb_r5;
    wire __A02_1__ovfstb_r6;
    wire __A02_2__EDSET;
    wire __A02_2__F01A;
    wire __A02_2__F01B;
    wire __A02_2__F01C;
    wire __A02_2__F01D;
    wire __A02_2__FS01;
    wire __A02_2__SB0;
    wire __A02_2__SB0_n;
    wire __A02_2__SB1;
    wire __A02_2__SB1_n;
    wire __A02_2__SB2;
    wire __A02_2__SB4;
    wire __A02_2__T12DC_n;
    wire __A02_2__TIMR;
    wire __A02_3__OVF;
    wire __A02_3__T01DC_n;
    wire __A02_3__T02DC_n;
    wire __A02_3__T03DC_n;
    wire __A02_3__T04DC_n;
    wire __A02_3__T05DC_n;
    wire __A02_3__T06DC_n;
    wire __A02_3__T07DC_n;
    wire __A02_3__T08DC_n;
    wire __A02_3__T09DC_n;
    wire __A02_3__T10DC_n;
    wand __A02_3__T12SET;
    wire __A02_3__T12SET_U2039_2;
    wire __A02_3__T12SET_U2039_4;
    wire __A02_3__T12SET_U2039_6;
    wire __A02_3__T12SET_U2039_8;
    wire __A02_3__UNF;
    wire __A02_NET_127;
    wire __A02_NET_141;
    wire __A02_NET_142;
    wire __A02_NET_143;
    wire __A02_NET_144;
    wire __A02_NET_145;
    wire __A02_NET_146;
    wire __A02_NET_147;
    wire __A02_NET_148;
    wire __A02_NET_149;
    wire __A02_NET_150;
    wire __A02_NET_151;
    wand __A02_NET_152;
    wire __A02_NET_152_U2020_2;
    wire __A02_NET_152_U2020_4;
    wire __A02_NET_153;
    wire __A02_NET_154;
    wire __A02_NET_155;
    wire __A02_NET_156;
    wire __A02_NET_157;
    wire __A02_NET_158;
    wire __A02_NET_159;
    wire __A02_NET_160;
    wire __A02_NET_161;
    wire __A02_NET_162;
    wire __A02_NET_163;
    wire __A02_NET_164;
    wire __A02_NET_165;
    wire __A02_NET_166;
    wire __A02_NET_167;
    wire __A02_NET_168;
    wire __A02_NET_169;
    wire __A02_NET_170;
    wire __A02_NET_171;
    wire __A02_NET_172;
    wire __A02_NET_173;
    wire __A02_NET_174;
    wire __A02_NET_175;
    wire __A02_NET_176;
    wire __A02_NET_177;
    wire __A02_NET_178;
    wire __A02_NET_179;
    wire __A02_NET_180;
    wire __A02_NET_181;
    wire __A02_NET_182;
    wire __A02_NET_183;
    wire __A02_NET_184;
    wire __A02_NET_185;
    wire __A02_NET_186;
    wire __A02_NET_187;
    wire __A02_NET_188;
    wire __A02_NET_189;
    wire __A02_NET_190;
    wire __A02_NET_191;
    wire __A02_NET_192;
    wire __A02_NET_193;
    wire __A02_NET_194;
    wire __A02_NET_195;
    wire __A02_NET_196;
    wire __A02_NET_197;
    wire __A02_NET_198;
    wire __A03_1__CSQG;
    wire __A03_1__IIP;
    wire __A03_1__IIP_n;
    wire __A03_1__INHINT;
    wire __A03_1__INKBT1;
    wire __A03_1__MIIP;
    wire __A03_1__MINHL;
    wire __A03_1__MSQ10;
    wire __A03_1__MSQ11;
    wire __A03_1__MSQ12;
    wire __A03_1__MSQ13;
    wire __A03_1__MSQ14;
    wire __A03_1__MSQ16;
    wire __A03_1__MSQEXT;
    wire __A03_1__NISQL;
    wire __A03_1__NISQL_n;
    wire __A03_1__QC0;
    wire __A03_1__RPTFRC;
    wire __A03_1__SQ3_n;
    wire __A03_1__SQ4_n;
    wire __A03_1__SQ5_n;
    wire __A03_1__SQ6_n;
    wire __A03_1__SQ7_n;
    wire __A03_1__SQEXT;
    wire __A03_1__SQR11;
    wire __A03_1__SQR12;
    wire __A03_1__SQR13;
    wire __A03_1__SQR14;
    wire __A03_1__SQR16;
    wire __A03_1__WSQG_n;
    wire __A03_1__wsqg;
    wire __A03_2__AUG0;
    wire __A03_2__BMF0;
    wire __A03_2__BMF0_n;
    wire __A03_2__BZF0;
    wire __A03_2__BZF0_n;
    wire __A03_2__DIM0;
    wand __A03_2__IC13_n;
    wire __A03_2__IC13_n_U3033_2;
    wire __A03_2__IC13_n_U3033_4;
    wire __A03_2__IC3_n;
    wire __A03_2__IC4_n;
    wire __A03_2__IC9_n;
    wire __A03_2__LXCH0;
    wire __A03_2__NDX0;
    wire __A03_2__NDXX1;
    wire __A03_2__NEXST0;
    wire __A03_2__NEXST0_n;
    wire __A03_2__QXCH0;
    wire __A03_2__SQ5QC0_n;
    wire __A03_2__TCSAJ3;
    wire __A03_NET_161;
    wire __A03_NET_163;
    wire __A03_NET_164;
    wire __A03_NET_165;
    wire __A03_NET_166;
    wire __A03_NET_167;
    wire __A03_NET_168;
    wire __A03_NET_169;
    wire __A03_NET_170;
    wire __A03_NET_171;
    wire __A03_NET_172;
    wire __A03_NET_174;
    wire __A03_NET_175;
    wire __A03_NET_176;
    wire __A03_NET_177;
    wire __A03_NET_178;
    wire __A03_NET_179;
    wire __A03_NET_180;
    wire __A03_NET_181;
    wire __A03_NET_182;
    wire __A03_NET_183;
    wire __A03_NET_184;
    wire __A03_NET_185;
    wire __A03_NET_186;
    wire __A03_NET_187;
    wire __A03_NET_188;
    wire __A03_NET_189;
    wire __A03_NET_190;
    wire __A03_NET_191;
    wire __A03_NET_192;
    wire __A03_NET_193;
    wire __A03_NET_194;
    wire __A03_NET_195;
    wire __A03_NET_196;
    wire __A03_NET_197;
    wire __A03_NET_198;
    wire __A03_NET_199;
    wire __A03_NET_200;
    wire __A03_NET_201;
    wire __A03_NET_202;
    wire __A03_NET_203;
    wire __A03_NET_204;
    wire __A03_NET_205;
    wire __A03_NET_206;
    wire __A03_NET_207;
    wire __A03_NET_208;
    wire __A03_NET_209;
    wire __A03_NET_210;
    wire __A03_NET_212;
    wire __A03_NET_213;
    wire __A03_NET_214;
    wire __A03_NET_215;
    wire __A03_NET_216;
    wire __A03_NET_217;
    wire __A03_NET_218;
    wire __A03_NET_219;
    wire __A03_NET_220;
    wire __A03_NET_221;
    wire __A03_NET_222;
    wire __A03_NET_223;
    wire __A03_NET_226;
    wire __A03_NET_227;
    wire __A03_NET_228;
    wire __A03_NET_229;
    wire __A03_NET_232;
    wire __A03_NET_233;
    wire __A04_1__DV0;
    wire __A04_1__DV0_n;
    wire __A04_1__DV376;
    wire __A04_1__DV3764;
    wire __A04_1__MBR1;
    wire __A04_1__MBR2;
    wire __A04_1__MST1;
    wire __A04_1__MST2;
    wire __A04_1__MST3;
    wand __A04_1__SGUM;
    wire __A04_1__SGUM_U4003_10;
    wire __A04_1__SGUM_U4003_12;
    wire __A04_1__ST1376_n;
    wire __A04_1__ST376;
    wire __A04_1__ST376_n;
    wire __A04_1__ST4_n;
    wire __A04_1__STG1;
    wire __A04_1__STG2;
    wire __A04_1__STG3;
    wire __A04_1__TSGN2;
    wire __A04_2__BR12B;
    wire __A04_2__BR1B2;
    wire __A04_2__BRXP3;
    wand __A04_2__L16_n;
    wire __A04_2__L16_n_U4063_8;
    wire __A04_2__MRSC;
    wire __A04_2__READ0_n;
    wire __A04_2__RUPT0_n;
    wire __A04_2__RUPT1_n;
    wire __A04_2__WOR0_n;
    wire __A04_2__WRITE0;
    wire __A04_2__WRITE0_n;
    wire __A04_NET_183;
    wire __A04_NET_184;
    wire __A04_NET_185;
    wire __A04_NET_186;
    wire __A04_NET_187;
    wire __A04_NET_188;
    wire __A04_NET_189;
    wire __A04_NET_190;
    wire __A04_NET_191;
    wire __A04_NET_192;
    wire __A04_NET_193;
    wire __A04_NET_194;
    wire __A04_NET_195;
    wire __A04_NET_196;
    wire __A04_NET_197;
    wire __A04_NET_198;
    wire __A04_NET_199;
    wire __A04_NET_200;
    wire __A04_NET_201;
    wire __A04_NET_202;
    wire __A04_NET_203;
    wire __A04_NET_204;
    wire __A04_NET_205;
    wire __A04_NET_206;
    wire __A04_NET_207;
    wire __A04_NET_210;
    wire __A04_NET_211;
    wand __A04_NET_212;
    wire __A04_NET_212_U4029_10;
    wire __A04_NET_212_U4029_8;
    wand __A04_NET_215;
    wire __A04_NET_215_U4023_6;
    wire __A04_NET_215_U4023_8;
    wand __A04_NET_216;
    wire __A04_NET_216_U4023_2;
    wire __A04_NET_216_U4023_4;
    wire __A04_NET_217;
    wire __A04_NET_218;
    wire __A04_NET_219;
    wire __A04_NET_220;
    wand __A04_NET_221;
    wire __A04_NET_221_U4023_10;
    wire __A04_NET_221_U4023_12;
    wire __A04_NET_221_U4029_2;
    wire __A04_NET_221_U4029_4;
    wire __A04_NET_221_U4029_6;
    wire __A04_NET_222;
    wire __A04_NET_223;
    wire __A04_NET_226;
    wire __A04_NET_227;
    wire __A04_NET_228;
    wire __A04_NET_229;
    wire __A04_NET_230;
    wire __A04_NET_231;
    wire __A04_NET_232;
    wire __A04_NET_233;
    wire __A04_NET_234;
    wire __A04_NET_235;
    wire __A04_NET_236;
    wire __A04_NET_237;
    wand __A04_NET_238;
    wire __A04_NET_238_U4003_6;
    wire __A04_NET_238_U4003_8;
    wire __A04_NET_239;
    wire __A04_NET_240;
    wire __A04_NET_241;
    wire __A04_NET_242;
    wire __A04_NET_243;
    wire __A04_NET_244;
    wire __A04_NET_245;
    wire __A04_NET_246;
    wire __A04_NET_247;
    wire __A04_NET_248;
    wire __A04_NET_249;
    wand __A04_NET_250;
    wire __A04_NET_250_U4003_2;
    wire __A04_NET_250_U4003_4;
    wire __A04_NET_251;
    wire __A04_NET_252;
    wire __A04_NET_253;
    wire __A04_NET_254;
    wire __A04_NET_255;
    wire __A04_NET_256;
    wire __A04_NET_259;
    wire __A04_NET_260;
    wire __A04_NET_261;
    wire __A04_NET_262;
    wire __A04_NET_263;
    wire __A04_NET_264;
    wire __A04_NET_265;
    wire __A04_NET_266;
    wire __A04_NET_267;
    wire __A04_NET_268;
    wire __A04_NET_269;
    wire __A04_NET_270;
    wire __A04_NET_271;
    wire __A04_NET_272;
    wire __A04_NET_273;
    wire __A04_NET_274;
    wire __A04_NET_275;
    wire __A04_NET_276;
    wire __A04_NET_277;
    wire __A04_NET_278;
    wire __A04_NET_279;
    wand __A04_NET_280;
    wire __A04_NET_280_U4045_4;
    wire __A04_NET_280_U4045_6;
    wire __A04_NET_281;
    wire __A04_NET_282;
    wire __A04_NET_283;
    wire __A04_NET_284;
    wire __A04_NET_285;
    wire __A04_NET_286;
    wire __A04_NET_287;
    wire __A04_NET_288;
    wire __A04_NET_289;
    wire __A04_NET_290;
    wire __A04_NET_291;
    wire __A04_NET_292;
    wire __A04_NET_293;
    wire __A04_NET_294;
    wire __A04_NET_295;
    wire __A04_NET_296;
    wire __A04_NET_297;
    wire __A04_NET_298;
    wire __A04_NET_299;
    wire __A04_NET_300;
    wire __A04_NET_301;
    wire __A04_NET_303;
    wire __A04_NET_306;
    wire __A04_NET_307;
    wire __A04_NET_308;
    wire __A04_NET_309;
    wire __A04_NET_310;
    wire __A04_NET_311;
    wire __A04_NET_312;
    wire __A04_NET_313;
    wire __A04_NET_314;
    wire __A04_NET_315;
    wire __A04_NET_316;
    wire __A04_NET_317;
    wire __A04_NET_318;
    wire __A04_NET_319;
    wire __A04_NET_320;
    wire __A04_NET_321;
    wire __A04_NET_322;
    wire __A04_NET_323;
    wire __A04_NET_324;
    wire __A04_NET_325;
    wire __A04_NET_326;
    wire __A04_NET_327;
    wire __A04_NET_328;
    wire __A04_NET_329;
    wire __A04_NET_330;
    wire __A04_NET_331;
    wire __A04_NET_332;
    wire __A04_NET_335;
    wire __A04_NET_336;
    wire __A04_NET_337;
    wire __A05_1__10XP6;
    wire __A05_1__10XP7;
    wire __A05_1__3XP5;
    wire __A05_1__8XP12;
    wire __A05_1__8XP15;
    wire __A05_1__8XP3;
    wire __A05_1__DV1B1B;
    wire __A05_1__GHNHC;
    wire __A05_1__MNISQ;
    wire __A05_1__NISQ_n;
    wire __A05_1__PARTC;
    wire __A05_1__PINC_n;
    wire __A05_1__RSTRT;
    wire __A05_2__10XP10;
    wire __A05_2__11XP6;
    wire __A05_2__5XP13;
    wire __A05_2__5XP19;
    wire __A05_2__5XP9;
    wire __A05_2__6XP2;
    wire __A05_2__6XP7;
    wire __A05_2__OCTAD3;
    wire __A05_2__OCTAD4;
    wire __A05_2__OCTAD5;
    wire __A05_2__OCTAD6;
    wire __A05_2__RSCT;
    wand __A05_2__Z15_n;
    wire __A05_2__Z15_n_U5067_2;
    wand __A05_2__Z16_n;
    wire __A05_2__Z16_n_U5058_4;
    wire __A05_NET_192;
    wire __A05_NET_194;
    wire __A05_NET_195;
    wire __A05_NET_196;
    wire __A05_NET_197;
    wire __A05_NET_198;
    wire __A05_NET_199;
    wire __A05_NET_200;
    wire __A05_NET_202;
    wire __A05_NET_203;
    wire __A05_NET_205;
    wire __A05_NET_206;
    wire __A05_NET_207;
    wire __A05_NET_208;
    wire __A05_NET_209;
    wire __A05_NET_210;
    wire __A05_NET_212;
    wire __A05_NET_213;
    wire __A05_NET_215;
    wire __A05_NET_216;
    wand __A05_NET_217;
    wire __A05_NET_217_U5035_2;
    wire __A05_NET_217_U5035_4;
    wire __A05_NET_217_U5035_6;
    wire __A05_NET_218;
    wire __A05_NET_219;
    wire __A05_NET_220;
    wire __A05_NET_221;
    wire __A05_NET_224;
    wire __A05_NET_225;
    wire __A05_NET_227;
    wire __A05_NET_228;
    wire __A05_NET_229;
    wire __A05_NET_230;
    wire __A05_NET_231;
    wire __A05_NET_232;
    wire __A05_NET_233;
    wire __A05_NET_234;
    wire __A05_NET_235;
    wire __A05_NET_236;
    wire __A05_NET_237;
    wire __A05_NET_238;
    wire __A05_NET_239;
    wire __A05_NET_240;
    wire __A05_NET_241;
    wire __A05_NET_242;
    wire __A05_NET_243;
    wire __A05_NET_244;
    wire __A05_NET_245;
    wire __A05_NET_246;
    wire __A05_NET_247;
    wire __A05_NET_248;
    wire __A05_NET_249;
    wire __A05_NET_250;
    wire __A05_NET_251;
    wire __A05_NET_252;
    wire __A05_NET_253;
    wire __A05_NET_254;
    wire __A05_NET_255;
    wire __A05_NET_256;
    wire __A05_NET_258;
    wire __A05_NET_259;
    wire __A05_NET_260;
    wire __A05_NET_261;
    wire __A05_NET_262;
    wire __A05_NET_263;
    wire __A05_NET_264;
    wire __A05_NET_265;
    wire __A05_NET_266;
    wire __A05_NET_267;
    wire __A05_NET_268;
    wire __A05_NET_269;
    wire __A05_NET_270;
    wire __A05_NET_271;
    wire __A05_NET_272;
    wire __A05_NET_273;
    wire __A05_NET_274;
    wire __A05_NET_275;
    wire __A05_NET_276;
    wire __A05_NET_277;
    wire __A05_NET_278;
    wire __A05_NET_279;
    wire __A05_NET_280;
    wire __A05_NET_281;
    wire __A05_NET_282;
    wire __A05_NET_283;
    wire __A05_NET_284;
    wire __A05_NET_285;
    wire __A05_NET_286;
    wire __A05_NET_287;
    wire __A05_NET_288;
    wire __A05_NET_289;
    wire __A05_NET_290;
    wire __A05_NET_291;
    wire __A05_NET_292;
    wire __A05_NET_294;
    wire __A05_NET_295;
    wire __A05_NET_296;
    wire __A05_NET_297;
    wire __A05_NET_298;
    wire __A05_NET_299;
    wire __A05_NET_300;
    wire __A05_NET_302;
    wire __A05_NET_303;
    wire __A05_NET_304;
    wire __A05_NET_305;
    wire __A05_NET_306;
    wire __A05_NET_308;
    wire __A05_NET_309;
    wire __A05_NET_310;
    wand __A05_NET_311;
    wire __A05_NET_311_U5035_10;
    wire __A05_NET_311_U5035_8;
    wire __A05_NET_312;
    wand __A05_NET_313;
    wire __A05_NET_313_U5041_6;
    wire __A05_NET_313_U5041_8;
    wire __A05_NET_314;
    wire __A05_NET_315;
    wire __A05_NET_316;
    wire __A05_NET_317;
    wire __A05_NET_318;
    wire __A05_NET_320;
    wire __A05_NET_321;
    wire __A05_NET_322;
    wire __A05_NET_323;
    wire __A05_NET_324;
    wire __A05_NET_326;
    wire __A05_NET_328;
    wire __A05_NET_329;
    wand __A05_NET_330;
    wire __A05_NET_330_U5051_12;
    wire __A05_NET_330_U5058_2;
    wire __A05_NET_331;
    wand __A05_NET_332;
    wire __A05_NET_332_U5058_10;
    wire __A05_NET_332_U5058_8;
    wire __A05_NET_333;
    wire __A05_NET_334;
    wire __A05_NET_335;
    wire __A05_NET_336;
    wire __A05_NET_338;
    wire __A05_NET_340;
    wire __A05_NET_342;
    wire __A05_NET_343;
    wire __A05_NET_344;
    wire __A05_NET_345;
    wire __A05_NET_346;
    wire __A05_NET_347;
    wire __A05_NET_348;
    wire __A05_NET_349;
    wire __A05_NET_350;
    wire __A05_NET_351;
    wire __A05_NET_352;
    wire __A05_NET_353;
    wire __A05_NET_354;
    wire __A05_NET_355;
    wire __A05_NET_356;
    wire __A05_NET_357;
    wire __A05_NET_358;
    wire __A05_NET_359;
    wire __A05_NET_360;
    wire __A05_NET_361;
    wire __A05_NET_362;
    wire __A05_NET_363;
    wire __A05_NET_364;
    wire __A05_NET_365;
    wire __A05_NET_366;
    wire __A05_NET_367;
    wire __A05_NET_368;
    wire __A05_NET_369;
    wire __A05_NET_370;
    wire __A05_NET_371;
    wire __A05_NET_372;
    wire __A05_NET_373;
    wire __A05_NET_374;
    wire __A06_1__DVXP1;
    wire __A06_1__L02A_n;
    wire __A06_1__L15A_n;
    wire __A06_1__RB1F;
    wire __A06_1__WHOMP_n;
    wire __A06_1__ZAP;
    wire __A06_1__ZIP;
    wire __A06_1__ZIPCI;
    wire __A06_2__10XP15;
    wire __A06_2__10XP9;
    wire __A06_2__6XP10;
    wire __A06_2__6XP12;
    wire __A06_2__7XP10;
    wire __A06_2__7XP11;
    wire __A06_2__7XP15;
    wire __A06_2__7XP7;
    wire __A06_2__8XP4;
    wire __A06_2__MOUT;
    wire __A06_2__POUT;
    wire __A06_2__PSEUDO;
    wire __A06_2__RDBANK;
    wire __A06_2__WOVR;
    wire __A06_2__ZOUT;
    wire __A06_NET_181;
    wire __A06_NET_182;
    wire __A06_NET_184;
    wire __A06_NET_185;
    wire __A06_NET_186;
    wire __A06_NET_187;
    wire __A06_NET_188;
    wire __A06_NET_189;
    wire __A06_NET_190;
    wire __A06_NET_191;
    wire __A06_NET_192;
    wire __A06_NET_193;
    wire __A06_NET_194;
    wire __A06_NET_195;
    wire __A06_NET_196;
    wire __A06_NET_199;
    wire __A06_NET_200;
    wire __A06_NET_201;
    wire __A06_NET_202;
    wand __A06_NET_203;
    wire __A06_NET_203_U6041_4;
    wire __A06_NET_203_U6041_6;
    wire __A06_NET_204;
    wire __A06_NET_205;
    wand __A06_NET_206;
    wire __A06_NET_206_U6041_10;
    wire __A06_NET_206_U6041_12;
    wire __A06_NET_207;
    wire __A06_NET_209;
    wire __A06_NET_210;
    wire __A06_NET_211;
    wire __A06_NET_212;
    wire __A06_NET_213;
    wire __A06_NET_216;
    wand __A06_NET_217;
    wire __A06_NET_217_U6019_10;
    wire __A06_NET_217_U6019_12;
    wire __A06_NET_218;
    wire __A06_NET_219;
    wire __A06_NET_220;
    wire __A06_NET_221;
    wire __A06_NET_222;
    wand __A06_NET_223;
    wire __A06_NET_223_U6029_2;
    wire __A06_NET_223_U6029_4;
    wire __A06_NET_224;
    wire __A06_NET_225;
    wire __A06_NET_229;
    wire __A06_NET_230;
    wire __A06_NET_232;
    wire __A06_NET_233;
    wire __A06_NET_234;
    wire __A06_NET_235;
    wire __A06_NET_237;
    wire __A06_NET_239;
    wire __A06_NET_240;
    wire __A06_NET_241;
    wire __A06_NET_242;
    wand __A06_NET_243;
    wire __A06_NET_243_U6047_10;
    wire __A06_NET_243_U6047_8;
    wire __A06_NET_244;
    wire __A06_NET_245;
    wire __A06_NET_246;
    wire __A06_NET_247;
    wire __A06_NET_248;
    wire __A06_NET_249;
    wire __A06_NET_250;
    wire __A06_NET_251;
    wire __A06_NET_252;
    wire __A06_NET_253;
    wire __A06_NET_254;
    wire __A06_NET_256;
    wire __A06_NET_257;
    wire __A06_NET_258;
    wire __A06_NET_259;
    wire __A06_NET_260;
    wire __A06_NET_261;
    wire __A06_NET_262;
    wire __A06_NET_263;
    wire __A06_NET_264;
    wire __A06_NET_266;
    wire __A06_NET_267;
    wire __A06_NET_268;
    wire __A06_NET_269;
    wire __A06_NET_270;
    wire __A06_NET_271;
    wire __A06_NET_272;
    wire __A06_NET_273;
    wire __A06_NET_274;
    wire __A06_NET_275;
    wire __A06_NET_276;
    wire __A06_NET_277;
    wire __A06_NET_278;
    wire __A06_NET_279;
    wand __A06_NET_280;
    wire __A06_NET_280_U6014_2;
    wire __A06_NET_280_U6014_4;
    wire __A06_NET_281;
    wire __A06_NET_282;
    wire __A06_NET_283;
    wire __A06_NET_284;
    wire __A06_NET_285;
    wire __A06_NET_286;
    wand __A06_NET_287;
    wire __A06_NET_287_U6004_2;
    wire __A06_NET_287_U6004_4;
    wire __A06_NET_288;
    wire __A06_NET_289;
    wire __A06_NET_290;
    wire __A06_NET_291;
    wire __A06_NET_292;
    wire __A06_NET_293;
    wire __A06_NET_294;
    wire __A06_NET_297;
    wire __A06_NET_298;
    wire __A06_NET_299;
    wire __A06_NET_300;
    wire __A06_NET_301;
    wire __A06_NET_302;
    wire __A06_NET_303;
    wire __A06_NET_304;
    wire __A06_NET_305;
    wire __A06_NET_306;
    wire __A06_NET_307;
    wire __A06_NET_309;
    wire __A06_NET_310;
    wire __A06_NET_311;
    wire __A06_NET_312;
    wire __A06_NET_313;
    wire __A06_NET_314;
    wire __A06_NET_315;
    wire __A06_NET_316;
    wire __A06_NET_317;
    wire __A06_NET_318;
    wire __A06_NET_319;
    wire __A06_NET_320;
    wire __A06_NET_321;
    wire __A06_NET_322;
    wire __A06_NET_323;
    wire __A06_NET_324;
    wire __A06_NET_325;
    wire __A06_NET_326;
    wire __A06_NET_327;
    wire __A06_NET_328;
    wire __A06_NET_329;
    wire __A06_NET_330;
    wire __A06_NET_334;
    wire __A06_NET_335;
    wire __A06_NET_336;
    wire __A06_NET_338;
    wire __A06_NET_339;
    wire __A06_NET_340;
    wire __A06_NET_341;
    wire __A06_NET_342;
    wire __A06_NET_343;
    wire __A06_NET_344;
    wire __A06_NET_345;
    wire __A06_NET_346;
    wire __A07_1__CCHG_n;
    wire __A07_1__MWAG;
    wire __A07_1__MWBG;
    wire __A07_1__MWG;
    wire __A07_1__MWLG;
    wire __A07_1__MWQG;
    wire __A07_1__MWSG;
    wire __A07_1__MWYG;
    wire __A07_1__MWZG;
    wire __A07_1__P04A;
    wire __A07_1__PIPSAM_n;
    wire __A07_1__WALSG;
    wire __A07_1__WCHG_n;
    wire __A07_1__WGA_n;
    wire __A07_1__WGNORM;
    wire __A07_1__WSCG_n;
    wire __A07_2__CEBG;
    wire __A07_2__CFBG;
    wire __A07_2__CIFF;
    wire __A07_2__CINORM;
    wire __A07_2__G2LSG;
    wire __A07_2__MRAG;
    wire __A07_2__MRGG;
    wire __A07_2__MRLG;
    wire __A07_2__MRULOG;
    wire __A07_2__MWBBEG;
    wire __A07_2__MWEBG;
    wire __A07_2__MWFBG;
    wire __A07_2__RBBEG_n;
    wire __A07_2__RBBK;
    wire __A07_2__RCHG_n;
    wire __A07_2__REBG_n;
    wire __A07_2__RFBG_n;
    wire __A07_2__RSCG_n;
    wire __A07_2__RUSG_n;
    wire __A07_2__U2BBKG_n;
    wire __A07_2__WBBEG_n;
    wire __A07_2__WEBG_n;
    wire __A07_2__WFBG_n;
    wire __A07_NET_137;
    wire __A07_NET_138;
    wire __A07_NET_139;
    wire __A07_NET_140;
    wire __A07_NET_141;
    wire __A07_NET_142;
    wire __A07_NET_143;
    wire __A07_NET_144;
    wire __A07_NET_145;
    wire __A07_NET_148;
    wire __A07_NET_149;
    wire __A07_NET_151;
    wire __A07_NET_152;
    wire __A07_NET_153;
    wire __A07_NET_154;
    wire __A07_NET_155;
    wire __A07_NET_156;
    wire __A07_NET_157;
    wire __A07_NET_158;
    wire __A07_NET_159;
    wire __A07_NET_160;
    wire __A07_NET_161;
    wand __A07_NET_162;
    wire __A07_NET_162_U7007_2;
    wire __A07_NET_162_U7007_4;
    wire __A07_NET_163;
    wire __A07_NET_164;
    wire __A07_NET_165;
    wire __A07_NET_166;
    wire __A07_NET_167;
    wire __A07_NET_168;
    wire __A07_NET_169;
    wire __A07_NET_170;
    wire __A07_NET_171;
    wire __A07_NET_172;
    wire __A07_NET_173;
    wire __A07_NET_174;
    wire __A07_NET_175;
    wire __A07_NET_177;
    wire __A07_NET_178;
    wire __A07_NET_179;
    wire __A07_NET_180;
    wire __A07_NET_181;
    wire __A07_NET_182;
    wire __A07_NET_183;
    wire __A07_NET_184;
    wire __A07_NET_185;
    wire __A07_NET_186;
    wire __A07_NET_187;
    wire __A07_NET_188;
    wire __A07_NET_189;
    wire __A07_NET_190;
    wire __A07_NET_191;
    wire __A07_NET_196;
    wire __A07_NET_197;
    wire __A07_NET_198;
    wire __A07_NET_199;
    wire __A07_NET_200;
    wire __A07_NET_201;
    wire __A07_NET_202;
    wire __A07_NET_203;
    wire __A07_NET_204;
    wire __A07_NET_205;
    wire __A07_NET_206;
    wire __A07_NET_207;
    wire __A07_NET_208;
    wire __A07_NET_209;
    wire __A07_NET_210;
    wire __A07_NET_211;
    wire __A07_NET_213;
    wire __A07_NET_214;
    wire __A08_1__X1;
    wire __A08_1__X1_n;
    wire __A08_1__X2;
    wire __A08_1__X2_n;
    wire __A08_1__Y1;
    wire __A08_1__Y1_n;
    wire __A08_1__Y2;
    wire __A08_1__Y2_n;
    wire __A08_1___A1_n;
    wire __A08_1___A2_n;
    wire __A08_1___B1_n;
    wire __A08_1___B2_n;
    wire __A08_1___CI_INTERNAL;
    wand __A08_1___G2_n;
    wire __A08_1___G2_n_U8028_10;
    wire __A08_1___G2_n_U8028_12;
    wire __A08_1___GEM1;
    wire __A08_1___GEM2;
    wire __A08_1___MWL1;
    wire __A08_1___MWL2;
    wire __A08_1___Q1_n;
    wire __A08_1___Q2_n;
    wand __A08_1___RL1_n;
    wire __A08_1___RL1_n_U8007_10;
    wire __A08_1___RL1_n_U8007_12;
    wire __A08_1___RL1_n_U8007_4;
    wire __A08_1___RL1_n_U8013_4;
    wand __A08_1___RL2_n;
    wire __A08_1___RL2_n_U8013_10;
    wire __A08_1___RL2_n_U8028_2;
    wire __A08_1___RL2_n_U8028_6;
    wire __A08_1___RL2_n_U8028_8;
    wire __A08_1___RL_OUT_1;
    wire __A08_1___RL_OUT_2;
    wire __A08_1___SUMA1;
    wire __A08_1___SUMA2;
    wire __A08_1___SUMB1;
    wire __A08_1___SUMB2;
    wire __A08_1___WL1;
    wire __A08_1___WL2;
    wand __A08_1___Z1_n;
    wire __A08_1___Z1_n_U8007_8;
    wand __A08_1___Z2_n;
    wire __A08_1___Z2_n_U8028_4;
    wire __A08_2__X1;
    wire __A08_2__X1_n;
    wire __A08_2__X2;
    wire __A08_2__X2_n;
    wire __A08_2__Y1;
    wire __A08_2__Y1_n;
    wire __A08_2__Y2;
    wire __A08_2__Y2_n;
    wire __A08_2___A1_n;
    wire __A08_2___A2_n;
    wire __A08_2___B1_n;
    wire __A08_2___B2_n;
    wire __A08_2___CI_IN;
    wire __A08_2___CI_INTERNAL;
    wand __A08_2___CO_IN;
    wire __A08_2___CO_IN_U8007_2;
    wire __A08_2___CO_IN_U8013_2;
    wand __A08_2___G1_n;
    wire __A08_2___G1_n_U8050_6;
    wire __A08_2___G1_n_U8050_8;
    wand __A08_2___G2_n;
    wire __A08_2___G2_n_U8063_10;
    wire __A08_2___G2_n_U8063_12;
    wire __A08_2___GEM1;
    wire __A08_2___GEM2;
    wand __A08_2___L1_n;
    wire __A08_2___L1_n_U8041_6;
    wire __A08_2___MWL1;
    wire __A08_2___MWL2;
    wire __A08_2___Q1_n;
    wire __A08_2___Q2_n;
    wand __A08_2___RL1_n;
    wire __A08_2___RL1_n_U8041_10;
    wire __A08_2___RL1_n_U8041_12;
    wire __A08_2___RL1_n_U8041_4;
    wire __A08_2___RL1_n_U8050_4;
    wand __A08_2___RL2_n;
    wire __A08_2___RL2_n_U8050_10;
    wire __A08_2___RL2_n_U8063_2;
    wire __A08_2___RL2_n_U8063_6;
    wire __A08_2___RL2_n_U8063_8;
    wire __A08_2___RL_OUT_1;
    wire __A08_2___RL_OUT_2;
    wire __A08_2___SUMA1;
    wire __A08_2___SUMA2;
    wire __A08_2___SUMB1;
    wire __A08_2___SUMB2;
    wire __A08_2___WL1;
    wire __A08_2___WL2;
    wire __A08_2___XUY1;
    wire __A08_2___XUY2;
    wand __A08_2___Z1_n;
    wire __A08_2___Z1_n_U8041_8;
    wand __A08_2___Z2_n;
    wire __A08_2___Z2_n_U8063_4;
    wire __A08_NET_137;
    wire __A08_NET_138;
    wire __A08_NET_139;
    wire __A08_NET_140;
    wire __A08_NET_141;
    wire __A08_NET_142;
    wire __A08_NET_143;
    wire __A08_NET_144;
    wire __A08_NET_145;
    wire __A08_NET_146;
    wire __A08_NET_147;
    wire __A08_NET_148;
    wire __A08_NET_149;
    wire __A08_NET_152;
    wire __A08_NET_155;
    wire __A08_NET_156;
    wire __A08_NET_157;
    wire __A08_NET_158;
    wire __A08_NET_159;
    wire __A08_NET_160;
    wire __A08_NET_161;
    wire __A08_NET_162;
    wire __A08_NET_163;
    wire __A08_NET_164;
    wire __A08_NET_167;
    wire __A08_NET_168;
    wire __A08_NET_169;
    wire __A08_NET_170;
    wire __A08_NET_173;
    wire __A08_NET_174;
    wire __A08_NET_175;
    wire __A08_NET_176;
    wire __A08_NET_177;
    wire __A08_NET_178;
    wire __A08_NET_179;
    wire __A08_NET_180;
    wire __A08_NET_181;
    wire __A08_NET_182;
    wire __A08_NET_183;
    wire __A08_NET_184;
    wire __A08_NET_185;
    wire __A08_NET_186;
    wire __A08_NET_187;
    wire __A08_NET_188;
    wire __A08_NET_189;
    wire __A08_NET_190;
    wire __A08_NET_191;
    wire __A08_NET_192;
    wire __A08_NET_193;
    wire __A08_NET_194;
    wire __A08_NET_195;
    wire __A08_NET_196;
    wire __A08_NET_197;
    wire __A08_NET_198;
    wire __A08_NET_199;
    wire __A08_NET_200;
    wire __A08_NET_205;
    wire __A08_NET_206;
    wire __A08_NET_207;
    wire __A08_NET_209;
    wire __A08_NET_210;
    wire __A08_NET_211;
    wire __A08_NET_212;
    wire __A08_NET_213;
    wire __A08_NET_214;
    wire __A08_NET_215;
    wire __A08_NET_216;
    wire __A08_NET_217;
    wire __A08_NET_218;
    wire __A08_NET_219;
    wire __A08_NET_220;
    wire __A08_NET_221;
    wire __A08_NET_222;
    wire __A08_NET_223;
    wire __A08_NET_224;
    wire __A08_NET_225;
    wire __A08_NET_226;
    wire __A08_NET_227;
    wire __A08_NET_228;
    wire __A08_NET_229;
    wire __A08_NET_230;
    wire __A08_NET_231;
    wire __A08_NET_232;
    wire __A08_NET_233;
    wire __A08_NET_234;
    wire __A08_NET_235;
    wire __A08_NET_236;
    wire __A08_NET_237;
    wire __A08_NET_238;
    wire __A08_NET_239;
    wire __A08_NET_240;
    wire __A08_NET_241;
    wire __A08_NET_242;
    wire __A08_NET_245;
    wire __A08_NET_248;
    wire __A08_NET_249;
    wire __A08_NET_250;
    wire __A08_NET_251;
    wire __A08_NET_252;
    wire __A08_NET_253;
    wire __A08_NET_254;
    wire __A08_NET_255;
    wire __A08_NET_256;
    wire __A08_NET_257;
    wire __A08_NET_260;
    wire __A08_NET_261;
    wire __A08_NET_262;
    wire __A08_NET_263;
    wire __A08_NET_266;
    wire __A08_NET_267;
    wire __A08_NET_268;
    wire __A08_NET_269;
    wire __A08_NET_270;
    wire __A08_NET_271;
    wire __A08_NET_272;
    wire __A08_NET_273;
    wire __A08_NET_274;
    wire __A08_NET_275;
    wire __A08_NET_276;
    wire __A08_NET_277;
    wire __A08_NET_278;
    wire __A08_NET_279;
    wire __A08_NET_280;
    wire __A08_NET_281;
    wire __A08_NET_282;
    wire __A08_NET_283;
    wire __A08_NET_284;
    wire __A08_NET_285;
    wire __A08_NET_286;
    wire __A08_NET_287;
    wire __A08_NET_288;
    wire __A08_NET_289;
    wire __A08_NET_290;
    wire __A08_NET_291;
    wire __A08_NET_293;
    wire __A08_NET_294;
    wire __A08_NET_298;
    wire __A08_NET_299;
    wire __A08_NET_300;
    wire __A08_NET_302;
    wire __A08_NET_303;
    wire __A08_NET_304;
    wire __A08_NET_305;
    wire __A08_NET_306;
    wire __A08_NET_307;
    wire __A08_NET_308;
    wire __A08_NET_309;
    wire __A08_NET_310;
    wire __A08_NET_311;
    wire __A08_NET_312;
    wire __A08_NET_313;
    wire __A08_NET_314;
    wire __A08_NET_315;
    wire __A08_NET_316;
    wire __A08_NET_317;
    wire __A08_NET_318;
    wire __A08_NET_319;
    wire __A08_NET_320;
    wire __A08_NET_321;
    wire __A08_NET_322;
    wire __A09_1__X1;
    wire __A09_1__X1_n;
    wire __A09_1__X2;
    wire __A09_1__X2_n;
    wire __A09_1__Y1;
    wire __A09_1__Y1_n;
    wire __A09_1__Y2;
    wire __A09_1__Y2_n;
    wire __A09_1___A1_n;
    wire __A09_1___A2_n;
    wire __A09_1___B1_n;
    wire __A09_1___B2_n;
    wire __A09_1___CI_INTERNAL;
    wire __A09_1___GEM1;
    wire __A09_1___GEM2;
    wand __A09_1___L1_n;
    wire __A09_1___L1_n_U9007_6;
    wand __A09_1___L2_n;
    wire __A09_1___L2_n_U9013_12;
    wire __A09_1___MWL1;
    wire __A09_1___MWL2;
    wire __A09_1___Q1_n;
    wire __A09_1___Q2_n;
    wand __A09_1___RL1_n;
    wire __A09_1___RL1_n_U9007_10;
    wire __A09_1___RL1_n_U9007_12;
    wire __A09_1___RL1_n_U9007_4;
    wire __A09_1___RL1_n_U9013_4;
    wand __A09_1___RL2_n;
    wire __A09_1___RL2_n_U9013_10;
    wire __A09_1___RL2_n_U9028_2;
    wire __A09_1___RL2_n_U9028_6;
    wire __A09_1___RL2_n_U9028_8;
    wire __A09_1___RL_OUT_1;
    wire __A09_1___RL_OUT_2;
    wire __A09_1___SUMA1;
    wire __A09_1___SUMA2;
    wire __A09_1___SUMB1;
    wire __A09_1___SUMB2;
    wire __A09_1___WL1;
    wire __A09_1___WL2;
    wand __A09_1___Z1_n;
    wire __A09_1___Z1_n_U9007_8;
    wand __A09_1___Z2_n;
    wire __A09_1___Z2_n_U9028_4;
    wire __A09_2__X1;
    wire __A09_2__X1_n;
    wire __A09_2__X2;
    wire __A09_2__X2_n;
    wire __A09_2__Y1;
    wire __A09_2__Y1_n;
    wire __A09_2__Y2;
    wire __A09_2__Y2_n;
    wire __A09_2___A1_n;
    wire __A09_2___A2_n;
    wire __A09_2___B1_n;
    wire __A09_2___B2_n;
    wire __A09_2___CI_IN;
    wire __A09_2___CI_INTERNAL;
    wand __A09_2___CO_IN;
    wire __A09_2___CO_IN_U9007_2;
    wire __A09_2___CO_IN_U9013_2;
    wand __A09_2___G2_n;
    wire __A09_2___G2_n_U9063_10;
    wire __A09_2___G2_n_U9063_12;
    wire __A09_2___GEM1;
    wire __A09_2___GEM2;
    wand __A09_2___L1_n;
    wire __A09_2___L1_n_U9041_6;
    wire __A09_2___MWL1;
    wire __A09_2___MWL2;
    wire __A09_2___Q1_n;
    wire __A09_2___Q2_n;
    wand __A09_2___RL1_n;
    wire __A09_2___RL1_n_U9041_10;
    wire __A09_2___RL1_n_U9041_12;
    wire __A09_2___RL1_n_U9041_4;
    wire __A09_2___RL1_n_U9050_4;
    wand __A09_2___RL2_n;
    wire __A09_2___RL2_n_U9050_10;
    wire __A09_2___RL2_n_U9063_2;
    wire __A09_2___RL2_n_U9063_6;
    wire __A09_2___RL2_n_U9063_8;
    wire __A09_2___RL_OUT_1;
    wire __A09_2___RL_OUT_2;
    wire __A09_2___SUMA1;
    wire __A09_2___SUMA2;
    wire __A09_2___SUMB1;
    wire __A09_2___SUMB2;
    wire __A09_2___WL1;
    wire __A09_2___WL2;
    wire __A09_2___XUY1;
    wire __A09_2___XUY2;
    wand __A09_2___Z1_n;
    wire __A09_2___Z1_n_U9041_8;
    wand __A09_2___Z2_n;
    wire __A09_2___Z2_n_U9063_4;
    wire __A09_NET_130;
    wire __A09_NET_131;
    wire __A09_NET_132;
    wire __A09_NET_133;
    wire __A09_NET_134;
    wire __A09_NET_135;
    wire __A09_NET_136;
    wire __A09_NET_137;
    wire __A09_NET_138;
    wire __A09_NET_139;
    wire __A09_NET_140;
    wire __A09_NET_141;
    wire __A09_NET_142;
    wire __A09_NET_145;
    wire __A09_NET_148;
    wire __A09_NET_149;
    wire __A09_NET_150;
    wire __A09_NET_151;
    wire __A09_NET_152;
    wire __A09_NET_153;
    wire __A09_NET_154;
    wire __A09_NET_155;
    wire __A09_NET_156;
    wire __A09_NET_157;
    wire __A09_NET_160;
    wire __A09_NET_161;
    wire __A09_NET_162;
    wire __A09_NET_163;
    wire __A09_NET_166;
    wire __A09_NET_167;
    wire __A09_NET_168;
    wire __A09_NET_169;
    wire __A09_NET_170;
    wire __A09_NET_171;
    wire __A09_NET_172;
    wire __A09_NET_173;
    wire __A09_NET_174;
    wire __A09_NET_175;
    wire __A09_NET_176;
    wire __A09_NET_177;
    wire __A09_NET_178;
    wire __A09_NET_179;
    wire __A09_NET_180;
    wire __A09_NET_181;
    wire __A09_NET_182;
    wire __A09_NET_183;
    wire __A09_NET_184;
    wire __A09_NET_185;
    wire __A09_NET_186;
    wire __A09_NET_187;
    wire __A09_NET_188;
    wire __A09_NET_189;
    wire __A09_NET_190;
    wire __A09_NET_191;
    wire __A09_NET_192;
    wire __A09_NET_193;
    wire __A09_NET_198;
    wire __A09_NET_199;
    wire __A09_NET_200;
    wire __A09_NET_202;
    wire __A09_NET_203;
    wire __A09_NET_204;
    wire __A09_NET_205;
    wire __A09_NET_206;
    wire __A09_NET_207;
    wire __A09_NET_208;
    wire __A09_NET_209;
    wire __A09_NET_210;
    wire __A09_NET_211;
    wire __A09_NET_212;
    wire __A09_NET_213;
    wire __A09_NET_214;
    wire __A09_NET_215;
    wire __A09_NET_216;
    wire __A09_NET_217;
    wire __A09_NET_218;
    wire __A09_NET_219;
    wire __A09_NET_220;
    wire __A09_NET_221;
    wire __A09_NET_222;
    wire __A09_NET_223;
    wire __A09_NET_224;
    wire __A09_NET_225;
    wire __A09_NET_226;
    wire __A09_NET_227;
    wire __A09_NET_228;
    wire __A09_NET_229;
    wire __A09_NET_230;
    wire __A09_NET_231;
    wire __A09_NET_232;
    wire __A09_NET_233;
    wire __A09_NET_234;
    wire __A09_NET_235;
    wire __A09_NET_238;
    wire __A09_NET_241;
    wire __A09_NET_242;
    wire __A09_NET_243;
    wire __A09_NET_244;
    wire __A09_NET_245;
    wire __A09_NET_246;
    wire __A09_NET_247;
    wire __A09_NET_248;
    wire __A09_NET_249;
    wire __A09_NET_250;
    wire __A09_NET_253;
    wire __A09_NET_254;
    wire __A09_NET_255;
    wire __A09_NET_256;
    wire __A09_NET_259;
    wire __A09_NET_260;
    wire __A09_NET_261;
    wire __A09_NET_262;
    wire __A09_NET_263;
    wire __A09_NET_264;
    wire __A09_NET_265;
    wire __A09_NET_266;
    wire __A09_NET_267;
    wire __A09_NET_268;
    wire __A09_NET_269;
    wire __A09_NET_270;
    wire __A09_NET_271;
    wire __A09_NET_272;
    wire __A09_NET_273;
    wire __A09_NET_274;
    wire __A09_NET_275;
    wire __A09_NET_276;
    wire __A09_NET_277;
    wire __A09_NET_278;
    wire __A09_NET_279;
    wire __A09_NET_280;
    wire __A09_NET_281;
    wire __A09_NET_282;
    wire __A09_NET_283;
    wire __A09_NET_284;
    wire __A09_NET_286;
    wire __A09_NET_287;
    wire __A09_NET_291;
    wire __A09_NET_292;
    wire __A09_NET_293;
    wire __A09_NET_295;
    wire __A09_NET_296;
    wire __A09_NET_297;
    wire __A09_NET_298;
    wire __A09_NET_299;
    wire __A09_NET_300;
    wire __A09_NET_301;
    wire __A09_NET_302;
    wire __A09_NET_303;
    wire __A09_NET_304;
    wire __A09_NET_305;
    wire __A09_NET_306;
    wire __A09_NET_307;
    wire __A09_NET_308;
    wire __A09_NET_309;
    wire __A09_NET_310;
    wire __A09_NET_311;
    wire __A09_NET_312;
    wire __A09_NET_313;
    wire __A09_NET_314;
    wire __A09_NET_315;
    wire __A10_1__X1;
    wire __A10_1__X1_n;
    wire __A10_1__X2;
    wire __A10_1__X2_n;
    wire __A10_1__Y1;
    wire __A10_1__Y1_n;
    wire __A10_1__Y2;
    wire __A10_1__Y2_n;
    wire __A10_1___A1_n;
    wire __A10_1___A2_n;
    wire __A10_1___B1_n;
    wire __A10_1___B2_n;
    wire __A10_1___CI_INTERNAL;
    wire __A10_1___GEM1;
    wire __A10_1___GEM2;
    wand __A10_1___L1_n;
    wire __A10_1___L1_n_U10007_6;
    wand __A10_1___L2_n;
    wire __A10_1___L2_n_U10013_12;
    wire __A10_1___MWL1;
    wire __A10_1___MWL2;
    wire __A10_1___Q1_n;
    wire __A10_1___Q2_n;
    wand __A10_1___RL1_n;
    wire __A10_1___RL1_n_U10007_10;
    wire __A10_1___RL1_n_U10007_12;
    wire __A10_1___RL1_n_U10007_4;
    wire __A10_1___RL1_n_U10013_4;
    wand __A10_1___RL2_n;
    wire __A10_1___RL2_n_U10013_10;
    wire __A10_1___RL2_n_U10028_2;
    wire __A10_1___RL2_n_U10028_6;
    wire __A10_1___RL2_n_U10028_8;
    wire __A10_1___RL_OUT_1;
    wire __A10_1___RL_OUT_2;
    wire __A10_1___SUMA1;
    wire __A10_1___SUMA2;
    wire __A10_1___SUMB1;
    wire __A10_1___SUMB2;
    wire __A10_1___WL1;
    wire __A10_1___WL2;
    wand __A10_1___Z1_n;
    wire __A10_1___Z1_n_U10007_8;
    wand __A10_1___Z2_n;
    wire __A10_1___Z2_n_U10028_4;
    wire __A10_2__X1;
    wire __A10_2__X1_n;
    wire __A10_2__X2;
    wire __A10_2__X2_n;
    wire __A10_2__Y1;
    wire __A10_2__Y1_n;
    wire __A10_2__Y2;
    wire __A10_2__Y2_n;
    wire __A10_2___A1_n;
    wire __A10_2___A2_n;
    wire __A10_2___B1_n;
    wire __A10_2___B2_n;
    wire __A10_2___CI_IN;
    wire __A10_2___CI_INTERNAL;
    wand __A10_2___CO_IN;
    wire __A10_2___CO_IN_U10007_2;
    wire __A10_2___CO_IN_U10013_2;
    wand __A10_2___G2_n;
    wire __A10_2___G2_n_U10063_10;
    wire __A10_2___G2_n_U10063_12;
    wire __A10_2___GEM1;
    wire __A10_2___GEM2;
    wand __A10_2___L1_n;
    wire __A10_2___L1_n_U10041_6;
    wire __A10_2___MWL1;
    wire __A10_2___MWL2;
    wire __A10_2___Q1_n;
    wire __A10_2___Q2_n;
    wand __A10_2___RL1_n;
    wire __A10_2___RL1_n_U10041_10;
    wire __A10_2___RL1_n_U10041_12;
    wire __A10_2___RL1_n_U10041_4;
    wire __A10_2___RL1_n_U10050_4;
    wand __A10_2___RL2_n;
    wire __A10_2___RL2_n_U10050_10;
    wire __A10_2___RL2_n_U10063_2;
    wire __A10_2___RL2_n_U10063_6;
    wire __A10_2___RL2_n_U10063_8;
    wire __A10_2___RL_OUT_1;
    wire __A10_2___RL_OUT_2;
    wire __A10_2___SUMA1;
    wire __A10_2___SUMA2;
    wire __A10_2___SUMB1;
    wire __A10_2___SUMB2;
    wire __A10_2___WL1;
    wire __A10_2___WL2;
    wire __A10_2___XUY1;
    wire __A10_2___XUY2;
    wand __A10_2___Z1_n;
    wire __A10_2___Z1_n_U10041_8;
    wand __A10_2___Z2_n;
    wire __A10_2___Z2_n_U10063_4;
    wire __A10_NET_129;
    wire __A10_NET_130;
    wire __A10_NET_131;
    wire __A10_NET_132;
    wire __A10_NET_133;
    wire __A10_NET_134;
    wire __A10_NET_135;
    wire __A10_NET_136;
    wire __A10_NET_137;
    wire __A10_NET_138;
    wire __A10_NET_139;
    wire __A10_NET_140;
    wire __A10_NET_141;
    wire __A10_NET_144;
    wire __A10_NET_147;
    wire __A10_NET_148;
    wire __A10_NET_149;
    wire __A10_NET_150;
    wire __A10_NET_151;
    wire __A10_NET_152;
    wire __A10_NET_153;
    wire __A10_NET_154;
    wire __A10_NET_155;
    wire __A10_NET_156;
    wire __A10_NET_159;
    wire __A10_NET_160;
    wire __A10_NET_161;
    wire __A10_NET_162;
    wire __A10_NET_165;
    wire __A10_NET_166;
    wire __A10_NET_167;
    wire __A10_NET_168;
    wire __A10_NET_169;
    wire __A10_NET_170;
    wire __A10_NET_171;
    wire __A10_NET_172;
    wire __A10_NET_173;
    wire __A10_NET_174;
    wire __A10_NET_175;
    wire __A10_NET_176;
    wire __A10_NET_177;
    wire __A10_NET_178;
    wire __A10_NET_179;
    wire __A10_NET_180;
    wire __A10_NET_181;
    wire __A10_NET_182;
    wire __A10_NET_183;
    wire __A10_NET_184;
    wire __A10_NET_185;
    wire __A10_NET_186;
    wire __A10_NET_187;
    wire __A10_NET_188;
    wire __A10_NET_189;
    wire __A10_NET_190;
    wire __A10_NET_191;
    wire __A10_NET_192;
    wire __A10_NET_197;
    wire __A10_NET_198;
    wire __A10_NET_199;
    wire __A10_NET_201;
    wire __A10_NET_202;
    wire __A10_NET_203;
    wire __A10_NET_204;
    wire __A10_NET_205;
    wire __A10_NET_206;
    wire __A10_NET_207;
    wire __A10_NET_208;
    wire __A10_NET_209;
    wire __A10_NET_210;
    wire __A10_NET_211;
    wire __A10_NET_212;
    wire __A10_NET_213;
    wire __A10_NET_214;
    wire __A10_NET_215;
    wire __A10_NET_216;
    wire __A10_NET_217;
    wire __A10_NET_218;
    wire __A10_NET_219;
    wire __A10_NET_220;
    wire __A10_NET_221;
    wire __A10_NET_222;
    wire __A10_NET_223;
    wire __A10_NET_224;
    wire __A10_NET_225;
    wire __A10_NET_226;
    wire __A10_NET_227;
    wire __A10_NET_228;
    wire __A10_NET_229;
    wire __A10_NET_230;
    wire __A10_NET_231;
    wire __A10_NET_232;
    wire __A10_NET_233;
    wire __A10_NET_234;
    wire __A10_NET_237;
    wire __A10_NET_240;
    wire __A10_NET_241;
    wire __A10_NET_242;
    wire __A10_NET_243;
    wire __A10_NET_244;
    wire __A10_NET_245;
    wire __A10_NET_246;
    wire __A10_NET_247;
    wire __A10_NET_248;
    wire __A10_NET_249;
    wire __A10_NET_252;
    wire __A10_NET_253;
    wire __A10_NET_254;
    wire __A10_NET_255;
    wire __A10_NET_258;
    wire __A10_NET_259;
    wire __A10_NET_260;
    wire __A10_NET_261;
    wire __A10_NET_262;
    wire __A10_NET_263;
    wire __A10_NET_264;
    wire __A10_NET_265;
    wire __A10_NET_266;
    wire __A10_NET_267;
    wire __A10_NET_268;
    wire __A10_NET_269;
    wire __A10_NET_270;
    wire __A10_NET_271;
    wire __A10_NET_272;
    wire __A10_NET_273;
    wire __A10_NET_274;
    wire __A10_NET_275;
    wire __A10_NET_276;
    wire __A10_NET_277;
    wire __A10_NET_278;
    wire __A10_NET_279;
    wire __A10_NET_280;
    wire __A10_NET_281;
    wire __A10_NET_282;
    wire __A10_NET_283;
    wire __A10_NET_285;
    wire __A10_NET_286;
    wire __A10_NET_290;
    wire __A10_NET_291;
    wire __A10_NET_292;
    wire __A10_NET_294;
    wire __A10_NET_295;
    wire __A10_NET_296;
    wire __A10_NET_297;
    wire __A10_NET_298;
    wire __A10_NET_299;
    wire __A10_NET_300;
    wire __A10_NET_301;
    wire __A10_NET_302;
    wire __A10_NET_303;
    wire __A10_NET_304;
    wire __A10_NET_305;
    wire __A10_NET_306;
    wire __A10_NET_307;
    wire __A10_NET_308;
    wire __A10_NET_309;
    wire __A10_NET_310;
    wire __A10_NET_311;
    wire __A10_NET_312;
    wire __A10_NET_313;
    wire __A10_NET_314;
    wire __A11_1__X1;
    wire __A11_1__X1_n;
    wire __A11_1__X2;
    wire __A11_1__X2_n;
    wire __A11_1__Y1;
    wire __A11_1__Y1_n;
    wire __A11_1__Y2;
    wire __A11_1__Y2_n;
    wire __A11_1___A1_n;
    wire __A11_1___A2_n;
    wire __A11_1___B1_n;
    wire __A11_1___B2_n;
    wire __A11_1___CI_INTERNAL;
    wire __A11_1___GEM1;
    wire __A11_1___GEM2;
    wand __A11_1___L1_n;
    wire __A11_1___L1_n_U11007_6;
    wand __A11_1___L2_n;
    wire __A11_1___L2_n_U11013_12;
    wire __A11_1___MWL1;
    wire __A11_1___MWL2;
    wire __A11_1___Q1_n;
    wire __A11_1___Q2_n;
    wand __A11_1___RL1_n;
    wire __A11_1___RL1_n_U11007_10;
    wire __A11_1___RL1_n_U11007_12;
    wire __A11_1___RL1_n_U11007_4;
    wire __A11_1___RL1_n_U11013_4;
    wand __A11_1___RL2_n;
    wire __A11_1___RL2_n_U11013_10;
    wire __A11_1___RL2_n_U11028_2;
    wire __A11_1___RL2_n_U11028_6;
    wire __A11_1___RL2_n_U11028_8;
    wire __A11_1___RL_OUT_1;
    wire __A11_1___RL_OUT_2;
    wire __A11_1___SUMA1;
    wire __A11_1___SUMA2;
    wire __A11_1___SUMB1;
    wire __A11_1___SUMB2;
    wire __A11_1___WL1;
    wire __A11_1___WL2;
    wand __A11_1___Z1_n;
    wire __A11_1___Z1_n_U11007_8;
    wand __A11_1___Z2_n;
    wire __A11_1___Z2_n_U11028_4;
    wire __A11_2__X1;
    wire __A11_2__X1_n;
    wire __A11_2__X2;
    wire __A11_2__X2_n;
    wire __A11_2__Y1;
    wire __A11_2__Y1_n;
    wire __A11_2__Y2;
    wire __A11_2__Y2_n;
    wire __A11_2___A1_n;
    wire __A11_2___A2_n;
    wire __A11_2___B1_n;
    wire __A11_2___B2_n;
    wire __A11_2___CI_IN;
    wire __A11_2___CI_INTERNAL;
    wand __A11_2___CO_IN;
    wire __A11_2___CO_IN_U11007_2;
    wire __A11_2___CO_IN_U11013_2;
    wand __A11_2___CO_OUT;
    wire __A11_2___CO_OUT_U11041_2;
    wire __A11_2___CO_OUT_U11050_2;
    wand __A11_2___G2_n;
    wire __A11_2___G2_n_U11063_10;
    wire __A11_2___G2_n_U11063_12;
    wire __A11_2___GEM1;
    wire __A11_2___GEM2;
    wand __A11_2___L2_n;
    wire __A11_2___L2_n_U11050_12;
    wire __A11_2___MWL1;
    wire __A11_2___MWL2;
    wire __A11_2___Q1_n;
    wire __A11_2___Q2_n;
    wand __A11_2___RL1_n;
    wire __A11_2___RL1_n_U11041_10;
    wire __A11_2___RL1_n_U11041_12;
    wire __A11_2___RL1_n_U11041_4;
    wire __A11_2___RL1_n_U11050_4;
    wand __A11_2___RL2_n;
    wire __A11_2___RL2_n_U11050_10;
    wire __A11_2___RL2_n_U11063_2;
    wire __A11_2___RL2_n_U11063_6;
    wire __A11_2___RL2_n_U11063_8;
    wire __A11_2___RL_OUT_1;
    wire __A11_2___RL_OUT_2;
    wire __A11_2___XUY1;
    wire __A11_2___XUY2;
    wand __A11_2___Z1_n;
    wire __A11_2___Z1_n_U11041_8;
    wand __A11_2___Z2_n;
    wire __A11_2___Z2_n_U11063_4;
    wire __A11_NET_130;
    wire __A11_NET_131;
    wire __A11_NET_132;
    wire __A11_NET_133;
    wire __A11_NET_134;
    wire __A11_NET_135;
    wire __A11_NET_136;
    wire __A11_NET_137;
    wire __A11_NET_138;
    wire __A11_NET_139;
    wire __A11_NET_140;
    wire __A11_NET_141;
    wire __A11_NET_142;
    wire __A11_NET_145;
    wire __A11_NET_148;
    wire __A11_NET_149;
    wire __A11_NET_150;
    wire __A11_NET_151;
    wire __A11_NET_152;
    wire __A11_NET_153;
    wire __A11_NET_154;
    wire __A11_NET_155;
    wire __A11_NET_156;
    wire __A11_NET_157;
    wire __A11_NET_160;
    wire __A11_NET_161;
    wire __A11_NET_162;
    wire __A11_NET_163;
    wire __A11_NET_166;
    wire __A11_NET_167;
    wire __A11_NET_168;
    wire __A11_NET_169;
    wire __A11_NET_170;
    wire __A11_NET_171;
    wire __A11_NET_172;
    wire __A11_NET_173;
    wire __A11_NET_174;
    wire __A11_NET_175;
    wire __A11_NET_176;
    wire __A11_NET_177;
    wire __A11_NET_178;
    wire __A11_NET_179;
    wire __A11_NET_180;
    wire __A11_NET_181;
    wire __A11_NET_182;
    wire __A11_NET_183;
    wire __A11_NET_184;
    wire __A11_NET_185;
    wire __A11_NET_186;
    wire __A11_NET_187;
    wire __A11_NET_188;
    wire __A11_NET_189;
    wire __A11_NET_190;
    wire __A11_NET_191;
    wire __A11_NET_192;
    wire __A11_NET_193;
    wire __A11_NET_198;
    wire __A11_NET_199;
    wire __A11_NET_200;
    wire __A11_NET_202;
    wire __A11_NET_203;
    wire __A11_NET_204;
    wire __A11_NET_205;
    wire __A11_NET_206;
    wire __A11_NET_207;
    wire __A11_NET_208;
    wire __A11_NET_209;
    wire __A11_NET_210;
    wire __A11_NET_211;
    wire __A11_NET_212;
    wire __A11_NET_213;
    wire __A11_NET_214;
    wire __A11_NET_215;
    wire __A11_NET_216;
    wire __A11_NET_217;
    wire __A11_NET_218;
    wire __A11_NET_219;
    wire __A11_NET_220;
    wire __A11_NET_221;
    wire __A11_NET_222;
    wire __A11_NET_223;
    wire __A11_NET_224;
    wire __A11_NET_225;
    wire __A11_NET_226;
    wire __A11_NET_227;
    wire __A11_NET_228;
    wire __A11_NET_229;
    wire __A11_NET_230;
    wire __A11_NET_231;
    wire __A11_NET_232;
    wire __A11_NET_233;
    wire __A11_NET_234;
    wire __A11_NET_235;
    wire __A11_NET_238;
    wire __A11_NET_241;
    wire __A11_NET_242;
    wire __A11_NET_243;
    wire __A11_NET_244;
    wire __A11_NET_245;
    wire __A11_NET_246;
    wire __A11_NET_247;
    wire __A11_NET_248;
    wire __A11_NET_249;
    wire __A11_NET_250;
    wire __A11_NET_253;
    wire __A11_NET_254;
    wire __A11_NET_255;
    wire __A11_NET_256;
    wire __A11_NET_259;
    wire __A11_NET_260;
    wire __A11_NET_261;
    wire __A11_NET_262;
    wire __A11_NET_263;
    wire __A11_NET_264;
    wire __A11_NET_265;
    wire __A11_NET_266;
    wire __A11_NET_267;
    wire __A11_NET_268;
    wire __A11_NET_269;
    wire __A11_NET_270;
    wire __A11_NET_271;
    wire __A11_NET_272;
    wire __A11_NET_273;
    wire __A11_NET_274;
    wire __A11_NET_275;
    wire __A11_NET_276;
    wire __A11_NET_277;
    wire __A11_NET_278;
    wire __A11_NET_279;
    wire __A11_NET_280;
    wire __A11_NET_281;
    wire __A11_NET_282;
    wire __A11_NET_283;
    wire __A11_NET_284;
    wire __A11_NET_286;
    wire __A11_NET_287;
    wire __A11_NET_291;
    wire __A11_NET_292;
    wire __A11_NET_293;
    wire __A11_NET_295;
    wire __A11_NET_296;
    wire __A11_NET_297;
    wire __A11_NET_298;
    wire __A11_NET_299;
    wire __A11_NET_300;
    wire __A11_NET_301;
    wire __A11_NET_302;
    wire __A11_NET_303;
    wire __A11_NET_304;
    wire __A11_NET_305;
    wire __A11_NET_306;
    wire __A11_NET_307;
    wire __A11_NET_308;
    wire __A11_NET_309;
    wire __A11_NET_310;
    wire __A11_NET_311;
    wire __A11_NET_312;
    wire __A11_NET_313;
    wire __A11_NET_314;
    wire __A11_NET_315;
    wire __A12_1__G01A_n;
    wire __A12_1__G02_n;
    wire __A12_1__G03_n;
    wire __A12_1__GEMP;
    wand __A12_1__GNZRO;
    wire __A12_1__GNZRO_U12016_2;
    wire __A12_1__GNZRO_U12016_4;
    wire __A12_1__MGP_n;
    wire __A12_1__MPAL;
    wire __A12_1__MSP;
    wire __A12_1__PA03;
    wire __A12_1__PA03_n;
    wire __A12_1__PA06;
    wire __A12_1__PA06_n;
    wire __A12_1__PA09;
    wire __A12_1__PA09_n;
    wire __A12_1__PA12;
    wire __A12_1__PA12_n;
    wire __A12_1__PA15;
    wire __A12_1__PA15_n;
    wand __A12_1__PALE;
    wire __A12_1__PALE_U12027_2;
    wire __A12_1__PALE_U12027_4;
    wire __A12_1__PB09;
    wire __A12_1__PB09_n;
    wire __A12_1__PB15;
    wire __A12_1__PB15_n;
    wire __A12_1__PC15;
    wire __A12_1__PC15_n;
    wire __A12_1__T7PHS4;
    wire __A12_1__T7PHS4_n;
    wire __A12_2__S01;
    wire __A12_2__S01_n;
    wire __A12_2__S02;
    wire __A12_2__S02_n;
    wire __A12_2__S03;
    wire __A12_2__S03_n;
    wire __A12_2__S04;
    wire __A12_2__S04_n;
    wire __A12_2__S05;
    wire __A12_2__S05_n;
    wire __A12_2__S06;
    wire __A12_2__S06_n;
    wire __A12_2__S07;
    wire __A12_2__S07_n;
    wire __A12_2__S08;
    wire __A12_2__S08_n;
    wire __A12_2__S09;
    wire __A12_2__S09_n;
    wire __A12_2__S10;
    wire __A12_2__S10_n;
    wire __A12_2__S11_n;
    wire __A12_2__S12_n;
    wire __A12_NET_106;
    wire __A12_NET_107;
    wire __A12_NET_108;
    wire __A12_NET_109;
    wire __A12_NET_110;
    wire __A12_NET_111;
    wire __A12_NET_112;
    wire __A12_NET_113;
    wire __A12_NET_114;
    wire __A12_NET_116;
    wire __A12_NET_118;
    wire __A12_NET_119;
    wire __A12_NET_120;
    wire __A12_NET_121;
    wire __A12_NET_122;
    wire __A12_NET_123;
    wire __A12_NET_124;
    wire __A12_NET_125;
    wire __A12_NET_126;
    wire __A12_NET_127;
    wire __A12_NET_128;
    wire __A12_NET_129;
    wire __A12_NET_130;
    wire __A12_NET_131;
    wire __A12_NET_132;
    wire __A12_NET_133;
    wire __A12_NET_134;
    wire __A12_NET_135;
    wire __A12_NET_136;
    wire __A12_NET_137;
    wire __A12_NET_138;
    wire __A12_NET_139;
    wire __A12_NET_140;
    wire __A12_NET_141;
    wire __A12_NET_142;
    wire __A12_NET_143;
    wire __A12_NET_146;
    wire __A12_NET_147;
    wire __A12_NET_148;
    wire __A12_NET_149;
    wire __A12_NET_150;
    wire __A12_NET_151;
    wire __A12_NET_155;
    wire __A12_NET_156;
    wire __A12_NET_165;
    wire __A12_NET_166;
    wire __A12_NET_168;
    wire __A12_NET_172;
    wire __A12_NET_173;
    wire __A12_NET_174;
    wire __A12_NET_177;
    wire __A12_NET_178;
    wire __A12_NET_179;
    wire __A12_NET_180;
    wire __A12_NET_181;
    wire __A12_NET_182;
    wire __A12_NET_183;
    wire __A12_NET_184;
    wire __A12_NET_185;
    wire __A12_NET_186;
    wire __A12_NET_189;
    wire __A12_NET_190;
    wire __A12_NET_191;
    wire __A12_NET_192;
    wire __A12_NET_193;
    wire __A12_NET_194;
    wire __A12_NET_195;
    wire __A12_NET_196;
    wire __A12_NET_197;
    wire __A12_NET_198;
    wire __A12_NET_199;
    wire __A12_NET_200;
    wire __A12_NET_204;
    wire __A12_NET_205;
    wire __A12_NET_206;
    wire __A12_NET_207;
    wire __A12_NET_208;
    wire __A12_NET_209;
    wire __A12_NET_210;
    wire __A12_NET_211;
    wire __A12_NET_212;
    wire __A12_NET_213;
    wire __A12_NET_214;
    wire __A12_NET_215;
    wire __A12_NET_216;
    wire __A12_NET_217;
    wire __A12_NET_218;
    wire __A12_NET_219;
    wire __A12_NET_220;
    wire __A12_NET_221;
    wire __A12_NET_222;
    wire __A12_NET_223;
    wire __A12_NET_224;
    wire __A12_NET_225;
    wire __A12_NET_226;
    wire __A12_NET_227;
    wire __A12_NET_228;
    wire __A12_NET_229;
    wire __A12_NET_230;
    wire __A12_NET_231;
    wire __A12_NET_232;
    wire __A12_NET_233;
    wire __A12_NET_234;
    wire __A12_NET_235;
    wire __A12_NET_236;
    wire __A12_NET_237;
    wire __A12_NET_238;
    wire __A12_NET_239;
    wire __A12_NET_240;
    wire __A12_NET_241;
    wire __A12_NET_242;
    wire __A12_NET_243;
    wire __A12_NET_244;
    wire __A12_NET_245;
    wire __A12_NET_246;
    wire __A12_NET_247;
    wire __A12_NET_248;
    wire __A12_NET_249;
    wire __A12_NET_250;
    wire __A12_NET_251;
    wire __A12_NET_252;
    wire n10XP1;
    wire n10XP8;
    wire n11XP2;
    wire n1XP10;
    wire n2XP3;
    wire n2XP5;
    wire n2XP7;
    wire n2XP8;
    wire n3XP2;
    wire n3XP6;
    wire n3XP7;
    wire n4XP11;
    wire n4XP5;
    wand n5XP11;
    wire n5XP11_U4039_6;
    wire n5XP11_U4039_8;
    wire n5XP12;
    wire n5XP15;
    wire n5XP21;
    wire n5XP28;
    wire n5XP4;
    wire n6XP5;
    wire n6XP8;
    wire n7XP14;
    wire n7XP19;
    wire n7XP4;
    wire n7XP9;
    wand n8PP4;
    wire n8PP4_U4063_12;
    wire n8PP4_U6037_10;
    wire n8PP4_U6037_12;
    wire n8PP4_U6041_2;
    wire n8XP5;
    wire n8XP6;
    wire n9XP1;
    wire n9XP5;



    U74HC02 #(1, 0, 1, 0) U1001(__A01_1__F02A, __A01_1__scaler_s2__FS_n, __A01_NET_169, __A01_1__F02B, __A01_NET_168, __A01_1__FS02, GND, __A01_NET_169, __A01_1__FS02, __A01_1__scaler_s2__FS_n, __A01_1__scaler_s2__FS_n, __A01_NET_168, __A01_1__FS02, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1002(__A01_1__F02A, FS01_n, __A01_NET_169, FS01_n, __A01_1__F02B, __A01_NET_168, GND, __A01_NET_171, __A01_1__F03A, __A01_1__F02A, __A01_NET_170, __A01_NET_169, __A01_NET_168, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1003(__A01_1__F03A, __A01_1__scaler_s3__FS_n, __A01_NET_171, __A01_1__F03B, __A01_NET_170, __A01_1__FS03, GND, __A01_NET_171, __A01_1__FS03, __A01_1__scaler_s3__FS_n, __A01_1__scaler_s3__FS_n, __A01_NET_170, __A01_1__FS03, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1004(__A01_NET_171, __A01_1__F02A, __A01_1__F04A, __A01_1__F03A, __A01_NET_172, __A01_NET_173, GND, __A01_NET_172, __A01_NET_173, __A01_1__F03A, __A01_1__F04B, __A01_NET_170, __A01_1__F03B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1005(__A01_1__F04A, __A01_1__scaler_s4__FS_n, __A01_NET_173, __A01_1__F04B, __A01_NET_172, __A01_1__FS04, GND, __A01_NET_173, __A01_1__FS04, __A01_1__scaler_s4__FS_n, __A01_1__scaler_s4__FS_n, __A01_NET_172, __A01_1__FS04, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1006(__A01_1__F05A, __A01_1__scaler_s5__FS_n, __A01_NET_174, __A01_1__F05B, __A01_NET_175, __A01_1__FS05, GND, __A01_NET_174, __A01_1__FS05, __A01_1__scaler_s5__FS_n, __A01_1__scaler_s5__FS_n, __A01_NET_175, __A01_1__FS05, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1007(__A01_1__F05A, __A01_1__F04A, __A01_NET_174, __A01_1__F04A, __A01_1__F05B, __A01_NET_175, GND, __A01_NET_176, __A01_1__F06A, __A01_1__F05A, __A01_NET_177, __A01_NET_174, __A01_NET_175, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1008(__A01_1__F06A, __A01_1__scaler_s6__FS_n, __A01_NET_176, __A01_1__F06B, __A01_NET_177, __A01_1__FS06, GND, __A01_NET_176, __A01_1__FS06, __A01_1__scaler_s6__FS_n, __A01_1__scaler_s6__FS_n, __A01_NET_177, __A01_1__FS06, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1009(__A01_NET_176, __A01_1__F05A, __A01_1__F07A, __A01_1__F06A, __A01_NET_178, __A01_NET_179, GND, __A01_NET_178, __A01_NET_179, __A01_1__F06A, __A01_1__F07B, __A01_NET_177, __A01_1__F06B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1010(__A01_1__F07A, __A01_1__scaler_s7__FS_n, __A01_NET_179, __A01_1__F07B, __A01_NET_178, __A01_1__FS07, GND, __A01_NET_179, __A01_1__FS07, __A01_1__scaler_s7__FS_n, __A01_1__scaler_s7__FS_n, __A01_NET_178, __A01_1__FS07, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1011(__A01_1__F08A, __A01_1__scaler_s8__FS_n, __A01_NET_181, __A01_1__F08B, __A01_NET_180, __A01_1__FS08, GND, __A01_NET_181, __A01_1__FS08, __A01_1__scaler_s8__FS_n, __A01_1__scaler_s8__FS_n, __A01_NET_180, __A01_1__FS08, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1012(__A01_1__F08A, __A01_1__F07A, __A01_NET_181, __A01_1__F07A, __A01_1__F08B, __A01_NET_180, GND, __A01_NET_183, __A01_1__F09A, __A01_1__F08A, __A01_NET_182, __A01_NET_181, __A01_NET_180, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1013(__A01_1__F09A, __A01_1__scaler_s9__FS_n, __A01_NET_183, __A01_1__F09B, __A01_NET_182, __A01_1__FS09, GND, __A01_NET_183, __A01_1__FS09, __A01_1__scaler_s9__FS_n, __A01_1__scaler_s9__FS_n, __A01_NET_182, __A01_1__FS09, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1014(__A01_NET_183, __A01_1__F08A, __A01_1__F10A, __A01_1__F09A, __A01_NET_184, __A01_NET_185, GND, __A01_NET_184, __A01_NET_185, __A01_1__F09A, __A01_1__F10B, __A01_NET_182, __A01_1__F09B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1015(__A01_1__F10A, __A01_1__scaler_s10__FS_n, __A01_NET_185, __A01_1__F10B, __A01_NET_184, __A01_1__FS10, GND, __A01_NET_185, __A01_1__FS10, __A01_1__scaler_s10__FS_n, __A01_1__scaler_s10__FS_n, __A01_NET_184, __A01_1__FS10, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1016(__A01_1__F11A, __A01_1__scaler_s11__FS_n, __A01_NET_187, __A01_1__F11B, __A01_NET_186, __A01_1__FS11, GND, __A01_NET_187, __A01_1__FS11, __A01_1__scaler_s11__FS_n, __A01_1__scaler_s11__FS_n, __A01_NET_186, __A01_1__FS11, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1017(__A01_1__F11A, __A01_1__F10A, __A01_NET_187, __A01_1__F10A, __A01_1__F11B, __A01_NET_186, GND, __A01_NET_188, __A01_1__F12A, __A01_1__F11A, __A01_NET_189, __A01_NET_187, __A01_NET_186, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1018(__A01_1__F12A, __A01_1__scaler_s12__FS_n, __A01_NET_188, __A01_1__F12B, __A01_NET_189, __A01_1__FS12, GND, __A01_NET_188, __A01_1__FS12, __A01_1__scaler_s12__FS_n, __A01_1__scaler_s12__FS_n, __A01_NET_189, __A01_1__FS12, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1019(__A01_NET_188, __A01_1__F11A, __A01_1__F13A, __A01_1__F12A, __A01_NET_190, __A01_NET_191, GND, __A01_NET_190, __A01_NET_191, __A01_1__F12A, __A01_1__F13B, __A01_NET_189, __A01_1__F12B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1020(__A01_1__F13A, __A01_1__scaler_s13__FS_n, __A01_NET_191, __A01_1__F13B, __A01_NET_190, __A01_1__FS13, GND, __A01_NET_191, __A01_1__FS13, __A01_1__scaler_s13__FS_n, __A01_1__scaler_s13__FS_n, __A01_NET_190, __A01_1__FS13, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1021(__A01_1__F14A, __A01_1__scaler_s14__FS_n, __A01_NET_193, __A01_1__F14B, __A01_NET_192, __A01_1__FS14, GND, __A01_NET_193, __A01_1__FS14, __A01_1__scaler_s14__FS_n, __A01_1__scaler_s14__FS_n, __A01_NET_192, __A01_1__FS14, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1022(__A01_1__F14A, __A01_1__F13A, __A01_NET_193, __A01_1__F13A, __A01_1__F14B, __A01_NET_192, GND, __A01_NET_195, __A01_1__F15A, __A01_1__F14A, __A01_NET_194, __A01_NET_193, __A01_NET_192, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1023(__A01_1__F15A, __A01_1__scaler_s15__FS_n, __A01_NET_195, __A01_1__F15B, __A01_NET_194, __A01_1__FS15, GND, __A01_NET_195, __A01_1__FS15, __A01_1__scaler_s15__FS_n, __A01_1__scaler_s15__FS_n, __A01_NET_194, __A01_1__FS15, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1024(__A01_NET_195, __A01_1__F14A, __A01_1__F16A, __A01_1__F15A, __A01_NET_197, __A01_NET_196, GND, __A01_NET_197, __A01_NET_196, __A01_1__F15A, __A01_1__F16B, __A01_NET_194, __A01_1__F15B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1025(__A01_1__F16A, __A01_1__scaler_s16__FS_n, __A01_NET_196, __A01_1__F16B, __A01_NET_197, __A01_1__FS16, GND, __A01_NET_196, __A01_1__FS16, __A01_1__scaler_s16__FS_n, __A01_1__scaler_s16__FS_n, __A01_NET_197, __A01_1__FS16, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1026(__A01_1__F17A, __A01_1__scaler_s17__FS_n, __A01_NET_199, __A01_1__F17B, __A01_NET_198, __A01_1__FS17, GND, __A01_NET_199, __A01_1__FS17, __A01_1__scaler_s17__FS_n, __A01_1__scaler_s17__FS_n, __A01_NET_198, __A01_1__FS17, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1027(__A01_1__F17A, __A01_1__F16A, __A01_NET_199, __A01_1__F16A, __A01_1__F17B, __A01_NET_198, GND,  ,  ,  ,  , __A01_NET_199, __A01_NET_198, VCC, SIM_RST, SIM_CLK);
    U74HC04 U1028(__A01_1__scaler_s2__FS_n, __A01_1__FS02A, __A01_1__scaler_s3__FS_n, __A01_1__FS03A, __A01_1__scaler_s4__FS_n, __A01_1__FS04A, GND, __A01_1__FS05A, __A01_1__scaler_s5__FS_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U1029(__A01_1__CHAT01, RCHAT_n, __A01_1__scaler_s6__FS_n, __A01_1__CHAT02, RCHAT_n, __A01_1__scaler_s7__FS_n, GND, RCHAT_n, __A01_1__scaler_s8__FS_n, __A01_1__CHAT03, RCHAT_n, __A01_1__scaler_s9__FS_n, __A01_1__CHAT04, VCC, SIM_RST, SIM_CLK);
    U74HC02 U1030(__A01_1__CHAT05, RCHAT_n, __A01_1__scaler_s10__FS_n, __A01_1__CHAT06, RCHAT_n, __A01_1__scaler_s11__FS_n, GND, RCHAT_n, __A01_1__scaler_s12__FS_n, __A01_1__CHAT07, RCHAT_n, __A01_1__scaler_s13__FS_n, __A01_1__CHAT08, VCC, SIM_RST, SIM_CLK);
    U74HC02 U1031(__A01_1__CHAT09, RCHAT_n, __A01_1__scaler_s14__FS_n, __A01_1__CHAT10, __A01_NET_143, __A01_1__scaler_s15__FS_n, GND, RCHAT_n, __A01_1__scaler_s16__FS_n, __A01_1__CHAT11, RCHAT_n, __A01_1__scaler_s17__FS_n, __A01_1__CHAT12, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1032(__A01_2__F18A, __A01_2__scaler_s18__FS_n, __A01_NET_201, __A01_2__F18B, __A01_NET_200, __A01_2__FS18, GND, __A01_NET_201, __A01_2__FS18, __A01_2__scaler_s18__FS_n, __A01_2__scaler_s18__FS_n, __A01_NET_200, __A01_2__FS18, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1033(__A01_2__F18A, __A01_1__F17A, __A01_NET_201, __A01_1__F17A, __A01_2__F18B, __A01_NET_200, GND, __A01_NET_203, __A01_2__F19A, __A01_2__F18A, __A01_NET_202, __A01_NET_201, __A01_NET_200, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1034(__A01_2__F19A, __A01_2__scaler_s19__FS_n, __A01_NET_203, __A01_2__F19B, __A01_NET_202, __A01_2__FS19, GND, __A01_NET_203, __A01_2__FS19, __A01_2__scaler_s19__FS_n, __A01_2__scaler_s19__FS_n, __A01_NET_202, __A01_2__FS19, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1035(__A01_NET_203, __A01_2__F18A, __A01_2__F20A, __A01_2__F19A, __A01_NET_204, __A01_NET_205, GND, __A01_NET_204, __A01_NET_205, __A01_2__F19A, __A01_2__F20B, __A01_NET_202, __A01_2__F19B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1036(__A01_2__F20A, __A01_2__scaler_s20__FS_n, __A01_NET_205, __A01_2__F20B, __A01_NET_204, __A01_2__FS20, GND, __A01_NET_205, __A01_2__FS20, __A01_2__scaler_s20__FS_n, __A01_2__scaler_s20__FS_n, __A01_NET_204, __A01_2__FS20, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1037(__A01_2__F21A, __A01_2__scaler_s21__FS_n, __A01_NET_207, __A01_2__F21B, __A01_NET_206, __A01_2__FS21, GND, __A01_NET_207, __A01_2__FS21, __A01_2__scaler_s21__FS_n, __A01_2__scaler_s21__FS_n, __A01_NET_206, __A01_2__FS21, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1038(__A01_2__F21A, __A01_2__F20A, __A01_NET_207, __A01_2__F20A, __A01_2__F21B, __A01_NET_206, GND, __A01_NET_209, __A01_2__F22A, __A01_2__F21A, __A01_NET_208, __A01_NET_207, __A01_NET_206, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1039(__A01_2__F22A, __A01_2__scaler_s22__FS_n, __A01_NET_209, __A01_2__F22B, __A01_NET_208, __A01_2__FS22, GND, __A01_NET_209, __A01_2__FS22, __A01_2__scaler_s22__FS_n, __A01_2__scaler_s22__FS_n, __A01_NET_208, __A01_2__FS22, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1040(__A01_NET_209, __A01_2__F21A, __A01_2__F23A, __A01_2__F22A, __A01_NET_210, __A01_NET_211, GND, __A01_NET_210, __A01_NET_211, __A01_2__F22A, __A01_2__F23B, __A01_NET_208, __A01_2__F22B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1041(__A01_2__F23A, __A01_2__scaler_s23__FS_n, __A01_NET_211, __A01_2__F23B, __A01_NET_210, __A01_2__FS23, GND, __A01_NET_211, __A01_2__FS23, __A01_2__scaler_s23__FS_n, __A01_2__scaler_s23__FS_n, __A01_NET_210, __A01_2__FS23, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1042(__A01_2__F24A, __A01_2__scaler_s24__FS_n, __A01_NET_213, __A01_2__F24B, __A01_NET_212, __A01_2__FS24, GND, __A01_NET_213, __A01_2__FS24, __A01_2__scaler_s24__FS_n, __A01_2__scaler_s24__FS_n, __A01_NET_212, __A01_2__FS24, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1043(__A01_2__F24A, __A01_2__F23A, __A01_NET_213, __A01_2__F23A, __A01_2__F24B, __A01_NET_212, GND, __A01_NET_215, __A01_2__F25A, __A01_2__F24A, __A01_NET_214, __A01_NET_213, __A01_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1044(__A01_2__F25A, __A01_2__scaler_s25__FS_n, __A01_NET_215, __A01_2__F25B, __A01_NET_214, __A01_2__FS25, GND, __A01_NET_215, __A01_2__FS25, __A01_2__scaler_s25__FS_n, __A01_2__scaler_s25__FS_n, __A01_NET_214, __A01_2__FS25, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1045(__A01_NET_215, __A01_2__F24A, __A01_2__F26A, __A01_2__F25A, __A01_NET_216, __A01_NET_217, GND, __A01_NET_216, __A01_NET_217, __A01_2__F25A, __A01_2__F26B, __A01_NET_214, __A01_2__F25B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1046(__A01_2__F26A, __A01_2__scaler_s26__FS_n, __A01_NET_217, __A01_2__F26B, __A01_NET_216, __A01_2__FS26, GND, __A01_NET_217, __A01_2__FS26, __A01_2__scaler_s26__FS_n, __A01_2__scaler_s26__FS_n, __A01_NET_216, __A01_2__FS26, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1047(__A01_2__F27A, __A01_2__scaler_s27__FS_n, __A01_NET_219, __A01_2__F27B, __A01_NET_218, __A01_2__FS27, GND, __A01_NET_219, __A01_2__FS27, __A01_2__scaler_s27__FS_n, __A01_2__scaler_s27__FS_n, __A01_NET_218, __A01_2__FS27, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1048(__A01_2__F27A, __A01_2__F26A, __A01_NET_219, __A01_2__F26A, __A01_2__F27B, __A01_NET_218, GND, __A01_NET_221, __A01_2__F28A, __A01_2__F27A, __A01_NET_220, __A01_NET_219, __A01_NET_218, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1049(__A01_2__F28A, __A01_2__scaler_s28__FS_n, __A01_NET_221, __A01_2__F28B, __A01_NET_220, __A01_2__FS28, GND, __A01_NET_221, __A01_2__FS28, __A01_2__scaler_s28__FS_n, __A01_2__scaler_s28__FS_n, __A01_NET_220, __A01_2__FS28, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1050(__A01_NET_221, __A01_2__F27A, __A01_2__F29A, __A01_2__F28A, __A01_NET_222, __A01_NET_223, GND, __A01_NET_222, __A01_NET_223, __A01_2__F28A, __A01_2__F29B, __A01_NET_220, __A01_2__F28B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1051(__A01_2__F29A, __A01_2__scaler_s29__FS_n, __A01_NET_223, __A01_2__F29B, __A01_NET_222, __A01_2__FS29, GND, __A01_NET_223, __A01_2__FS29, __A01_2__scaler_s29__FS_n, __A01_2__scaler_s29__FS_n, __A01_NET_222, __A01_2__FS29, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1052(__A01_2__F30A, __A01_2__scaler_s30__FS_n, __A01_NET_225, __A01_2__F30B, __A01_NET_224, __A01_2__FS30, GND, __A01_NET_225, __A01_2__FS30, __A01_2__scaler_s30__FS_n, __A01_2__scaler_s30__FS_n, __A01_NET_224, __A01_2__FS30, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1053(__A01_2__F30A, __A01_2__F29A, __A01_NET_225, __A01_2__F29A, __A01_2__F30B, __A01_NET_224, GND, __A01_NET_227, __A01_2__F31A, __A01_2__F30A, __A01_NET_226, __A01_NET_225, __A01_NET_224, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1054(__A01_2__F31A, __A01_2__scaler_s31__FS_n, __A01_NET_227, __A01_2__F31B, __A01_NET_226, __A01_2__FS31, GND, __A01_NET_227, __A01_2__FS31, __A01_2__scaler_s31__FS_n, __A01_2__scaler_s31__FS_n, __A01_NET_226, __A01_2__FS31, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1055(__A01_NET_227, __A01_2__F30A, __A01_2__F32A, __A01_2__F31A, __A01_NET_228, __A01_NET_229, GND, __A01_NET_228, __A01_NET_229, __A01_2__F31A, __A01_2__F32B, __A01_NET_226, __A01_2__F31B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1056(__A01_2__F32A, __A01_2__scaler_s32__FS_n, __A01_NET_229, __A01_2__F32B, __A01_NET_228, __A01_2__FS32, GND, __A01_NET_229, __A01_2__FS32, __A01_2__scaler_s32__FS_n, __A01_2__scaler_s32__FS_n, __A01_NET_228, __A01_2__FS32, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U1057(__A01_2__F33A, __A01_2__scaler_s33__FS_n, __A01_NET_231, __A01_2__F33B, __A01_NET_230, __A01_2__FS33, GND, __A01_NET_231, __A01_2__FS33, __A01_2__scaler_s33__FS_n, __A01_2__scaler_s33__FS_n, __A01_NET_230, __A01_2__FS33, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1058(__A01_2__F33A, __A01_2__F32A, __A01_NET_231, __A01_2__F32A, __A01_2__F33B, __A01_NET_230, GND,  ,  ,  ,  , __A01_NET_231, __A01_NET_230, VCC, SIM_RST, SIM_CLK);
    U74HC02 U1059(__A01_2__CHAT13, RCHAT_n, __A01_2__scaler_s18__FS_n, __A01_2__CHAT14, RCHAT_n, __A01_2__scaler_s19__FS_n, GND, RCHBT_n, __A01_2__scaler_s20__FS_n, __A01_2__CHBT01, RCHBT_n, __A01_2__scaler_s21__FS_n, __A01_2__CHBT02, VCC, SIM_RST, SIM_CLK);
    U74HC02 U1060(__A01_2__CHBT03, RCHBT_n, __A01_2__scaler_s22__FS_n, __A01_2__CHBT04, RCHBT_n, __A01_2__scaler_s23__FS_n, GND, RCHBT_n, __A01_2__scaler_s24__FS_n, __A01_2__CHBT05, RCHBT_n, __A01_2__scaler_s25__FS_n, __A01_2__CHBT06, VCC, SIM_RST, SIM_CLK);
    U74HC02 U1061(__A01_2__CHBT07, RCHBT_n, __A01_2__scaler_s26__FS_n, __A01_2__CHBT08, RCHBT_n, __A01_2__scaler_s27__FS_n, GND, RCHBT_n, __A01_2__scaler_s28__FS_n, __A01_2__CHBT09, RCHBT_n, __A01_2__scaler_s29__FS_n, __A01_2__CHBT10, VCC, SIM_RST, SIM_CLK);
    U74HC02 U1062(__A01_2__CHBT11, RCHBT_n, __A01_2__scaler_s30__FS_n, __A01_2__CHBT12, __A01_NET_155, __A01_2__scaler_s31__FS_n, GND, RCHBT_n, __A01_2__scaler_s32__FS_n, __A01_2__CHBT13, RCHBT_n, __A01_2__scaler_s33__FS_n, __A01_2__CHBT14, VCC, SIM_RST, SIM_CLK);


    U74HC02 #(0, 1, 0, 0) U2001(__A02_1__cdiv_1__D, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__B, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__B, __A02_1__cdiv_1__FS, GND, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__A, __A02_1__cdiv_1__FS, __A02_1__cdiv_1__A, __A02_1__cdiv_1__FS, PHS2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U2002(__A02_1__cdiv_1__D, CLOCK, __A02_1__cdiv_1__B, CLOCK, PHS2, __A02_1__cdiv_1__A, GND, __A02_2__EDSET, P02, P03_n, P04, __A02_1__cdiv_1__B, __A02_1__cdiv_1__A, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1, 0, 0, 1, 0, 1) U2003(__A02_1__cdiv_1__D, __A02_1__cdiv_2__F, PHS2, PHS2_n, PHS4, PHS4_n, GND, __A02_NET_127, __A02_1__cdiv_1__B, CT, __A02_NET_127, CT_n, CT, VCC, SIM_RST, SIM_CLK);
    U74HC02 U2004(PHS4, __A02_1__cdiv_2__F, __A02_1__cdiv_1__A, __A02_1__oddset, STOP, __A02_1__RINGA_n, GND, P02_n, P04, __A02_2__SB4, P01, __A02_NET_154, __A02_NET_155, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(0, 0, 0, 0, 1, 1) U2005(__A02_1__cdiv_1__FS_n, WT, WT, WT_n, WT, TT_n, GND, __A02_1__ovfstb_r5, __A02_1__ovfstb_r4, __A02_1__ovfstb_r6, __A02_1__ovfstb_r5, __A02_1__OVFSTB_n, __A02_1__ovfstb_r2, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U2006(__A02_1__cdiv_2__D, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__FS, GND, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__A, __A02_1__cdiv_2__FS, __A02_1__cdiv_2__A, __A02_1__cdiv_2__FS, __A02_1__cdiv_2__C, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U2007(__A02_1__cdiv_2__D, __A02_1__cdiv_2__F, __A02_1__cdiv_2__B, __A02_1__cdiv_2__F, __A02_1__cdiv_2__C, __A02_1__cdiv_2__A, GND, P03, __A02_2__EDSET, __A02_NET_168, P03_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__A, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1, 0, 1, 0, 0, 0) U2008(__A02_1__cdiv_2__D, __A02_1__RINGA_n, __A02_1__oddset, __A02_1__ODDSET_n, __A02_1__cdiv_2__C, __A02_1__RINGB_n, GND, __A02_1__evnset, __A02_1__RINGB_n, __A02_1__EVNSET_n, __A02_1__evnset, RT, __A02_1__cdiv_1__A, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 0, 1) U2009(__A02_1__ovfstb_r1, CT_n, __A02_1__ovfstb_r2, __A02_1__ovfstb_r2, __A02_1__ovfstb_r6, __A02_1__ovfstb_r1, GND, __A02_1__ovfstb_r4, __A02_1__ovfstb_r2, __A02_1__ovfstb_r3, __A02_1__ovfstb_r3, __A02_1__ovfstb_r1, __A02_1__ovfstb_r4, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1, 0, 0, 0, 0, 0) U2010(CT, PHS3_n, WT_n, CLK, WT_n, MONWT, GND, Q2A, WT_n, RT_n, RT, __A02_2__TIMR, __A02_NET_159, VCC, SIM_RST, SIM_CLK);
    U74HC27 U2011(__A02_1__RINGB_n, P05_n, P04, P05, __A02_1__RINGA_n, __A02_NET_166, GND, __A02_NET_148, __A02_2__T12DC_n, __A02_NET_152, __A02_1__EVNSET_n, __A02_NET_164, P04_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U2012(P01, __A02_NET_164, P01_n, P01_n, P01, __A02_NET_166, GND, __A02_1__RINGA_n, P01, __A02_NET_169, P01_n, __A02_1__RINGB_n, __A02_NET_167, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U2013(P02, __A02_NET_169, P02_n, P02_n, P02, __A02_NET_167, GND, __A02_1__RINGB_n, P02, __A02_NET_168, P02_n, __A02_1__RINGA_n, __A02_NET_162, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U2014(__A02_NET_154, __A02_NET_155, STOP_n, P03_n, P03, __A02_NET_162, GND, __A02_1__RINGA_n, P03, __A02_NET_161, P03_n, __A02_1__RINGB_n, __A02_NET_160, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U2015(P04, __A02_NET_161, P04_n, P04_n, P04, __A02_NET_160, GND, __A02_1__RINGB_n, P04, __A02_NET_165, P04_n, __A02_1__RINGA_n, __A02_NET_163, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U2016(P05, __A02_NET_165, P05_n, P05_n, P05, __A02_NET_163, GND, __A02_NET_152, GOJ1, __A02_NET_153, __A02_1__EVNSET_n, __A02_NET_147, __A02_NET_149, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U2017(__A02_2__F01D, FS01_n, __A02_2__F01B, FS01_n, __A02_2__F01B, __A02_2__FS01, GND, FS01_n, __A02_2__F01A, __A02_2__FS01, __A02_2__F01A, __A02_2__FS01, __A02_2__F01C, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U2018(__A02_2__F01D, P01_n, __A02_2__F01B, P01_n, __A02_2__F01C, __A02_2__F01A, GND,  ,  ,  ,  , __A02_2__F01B, __A02_2__F01A, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 1, 0) U2019(SBY, ALGA, STRT1, STRT2, __A02_NET_153, __A02_NET_151, GND, __A02_NET_146, __A02_2__T12DC_n, __A02_NET_141, __A02_1__EVNSET_n, __A02_NET_150, MSTRTP, VCC, SIM_RST, SIM_CLK);
    assign __A02_NET_152 = __A02_NET_152_U2020_2;
    assign __A02_NET_152 = __A02_NET_152_U2020_4;
    U74LVC07 U2020(__A02_NET_150, __A02_NET_152_U2020_2, __A02_NET_151, __A02_NET_152_U2020_4,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1, 0, 1, 0, 1, 0) U2021(__A02_NET_152, __A02_NET_147, MSTP, __A02_NET_141, GOJAM_n, GOJAM, GND, MGOJAM, GOJAM, STOP, STOP_n, MSTPIT_n, STOP, VCC, SIM_RST, SIM_CLK);
    U74HC02 U2022(__A02_NET_142, __A02_1__EVNSET_n, MSTP, GOJAM_n, STRT2, STOPA, GND, STOPA, __A02_NET_145, STOP_n, STRT2, __A02_NET_158, __A02_NET_159, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 1) U2023(__A02_NET_143, __A02_NET_148, STOPA, STOPA, __A02_NET_143, __A02_NET_149, GND, __A02_NET_146, __A02_NET_145, __A02_NET_144, __A02_NET_144, __A02_NET_142, __A02_NET_145, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U2024(__A02_3__T12SET, GOJAM, __A02_3__T01DC_n, __A02_NET_193, GOJAM, __A02_NET_190, GND, __A02_NET_193, __A02_3__T02DC_n, __A02_NET_192, GOJAM, __A02_2__T12DC_n, __A02_NET_191, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 0, 1) U2025(__A02_NET_191, __A02_2__T12DC_n, __A02_NET_190, __A02_NET_181, __A02_2__T12DC_n, __A02_1__ODDSET_n, GND, __A02_2__T12DC_n, __A02_1__EVNSET_n, T12, __A02_NET_181, __A02_NET_190, __A02_3__T01DC_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U2026(__A02_NET_180, __A02_3__T01DC_n, __A02_1__EVNSET_n, T01, __A02_3__T01DC_n, __A02_1__ODDSET_n, GND, __A02_NET_180, __A02_NET_193, __A02_3__T02DC_n, __A02_3__T02DC_n, __A02_1__ODDSET_n, __A02_NET_185, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U2027(T02, __A02_3__T02DC_n, __A02_1__EVNSET_n, __A02_3__T03DC_n, __A02_NET_185, __A02_NET_192, GND, __A02_3__T03DC_n, __A02_1__EVNSET_n, __A02_NET_186, __A02_3__T03DC_n, __A02_1__ODDSET_n, T03, VCC, SIM_RST, SIM_CLK);
    U74HC27 U2028(__A02_3__T03DC_n, __A02_NET_188, __A02_3__T04DC_n, __A02_NET_187, GOJAM, __A02_NET_188, GND, __A02_NET_187, __A02_3__T05DC_n, __A02_NET_189, GOJAM, __A02_NET_192, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 0, 1) U2029(__A02_3__T04DC_n, __A02_NET_186, __A02_NET_188, __A02_NET_183, __A02_3__T04DC_n, __A02_1__ODDSET_n, GND, __A02_3__T04DC_n, __A02_1__EVNSET_n, T04, __A02_NET_183, __A02_NET_187, __A02_3__T05DC_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U2030(__A02_NET_174, __A02_3__T05DC_n, __A02_1__EVNSET_n, T05, __A02_3__T05DC_n, __A02_1__ODDSET_n, GND, __A02_NET_189, __A02_NET_174, __A02_3__T06DC_n, __A02_1__EVNSET_n, __A02_3__T06DC_n, T06, VCC, SIM_RST, SIM_CLK);
    U74HC27 U2031(GOJAM, __A02_NET_196, GOJAM, __A02_NET_195, __A02_3__T07DC_n, __A02_NET_196, GND, __A02_NET_195, GOJAM, __A02_NET_198, __A02_3__T08DC_n, __A02_NET_189, __A02_3__T06DC_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U2032(__A02_NET_182, __A02_1__ODDSET_n, __A02_3__T06DC_n, __A02_3__T07DC_n, __A02_NET_196, __A02_NET_182, GND, __A02_1__ODDSET_n, __A02_3__T07DC_n, T07, __A02_1__EVNSET_n, __A02_3__T07DC_n, __A02_NET_184, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 0, 1) U2033(__A02_3__T08DC_n, __A02_NET_195, __A02_NET_184, T08, __A02_1__EVNSET_n, __A02_3__T08DC_n, GND, __A02_1__ODDSET_n, __A02_3__T08DC_n, __A02_NET_176, __A02_NET_198, __A02_NET_176, __A02_3__T09DC_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U2034(GOJAM, __A02_NET_197, GOJAM, __A02_NET_194, __A02_3__T10DC_n, __A02_NET_197, GND, __A02_NET_194, GOJAM, __A02_NET_177, __A02_NET_179, __A02_NET_198, __A02_3__T09DC_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U2035(T09, __A02_1__ODDSET_n, __A02_3__T09DC_n, __A02_NET_175, __A02_1__EVNSET_n, __A02_3__T09DC_n, GND, __A02_NET_197, __A02_NET_175, __A02_3__T10DC_n, __A02_1__EVNSET_n, __A02_NET_197, __A02_NET_177, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U2036(__A02_NET_178, __A02_1__ODDSET_n, __A02_3__T10DC_n, __A02_NET_179, __A02_NET_194, __A02_NET_178, GND, __A02_1__EVNSET_n, __A02_3__T10DC_n, T10, __A02_1__ODDSET_n, __A02_NET_179, T11, VCC, SIM_RST, SIM_CLK);
    U74HC02 U2037(__A02_NET_170, __A02_NET_193, __A02_NET_190, __A02_2__SB0, P02_n, P05, GND, P05_n, P03_n, __A02_2__SB1, P05_n, P02, __A02_2__SB2, VCC, SIM_RST, SIM_CLK);
    U74HC27 U2038(__A02_NET_187, __A02_NET_188, __A02_NET_198, __A02_NET_197, __A02_1__EVNSET_n, __A02_NET_172, GND, __A02_NET_173, __A02_NET_189, __A02_NET_196, __A02_NET_195, __A02_NET_171, __A02_NET_192, VCC, SIM_RST, SIM_CLK);
    assign __A02_3__T12SET = __A02_3__T12SET_U2039_2;
    assign __A02_3__T12SET = __A02_3__T12SET_U2039_4;
    assign __A02_3__T12SET = __A02_3__T12SET_U2039_6;
    assign __A02_3__T12SET = __A02_3__T12SET_U2039_8;
    U74LVC07 U2039(__A02_NET_170, __A02_3__T12SET_U2039_2, __A02_NET_171, __A02_3__T12SET_U2039_4, __A02_NET_172, __A02_3__T12SET_U2039_6, GND, __A02_3__T12SET_U2039_8, __A02_NET_173,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1, 0, 1, 0, 1, 0) U2040(T01, T01_n, T01_n, MT01, T02, T02_n, GND, MT02, T02_n, T03_n, T03, MT03, T03_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1, 0, 1, 0, 1, 0) U2041(T04, T04_n, T04_n, MT04, T05, T05_n, GND, MT05, T05_n, T06_n, T06, MT06, T06_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1, 0, 1, 0, 1, 0) U2042(T07, T07_n, T07_n, MT07, T08, T08_n, GND, MT08, T08_n, T09_n, T09, MT09, T09_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1, 0, 1, 0, 1, 0) U2043(T10, T10_n, T10_n, MT10, T11, T11_n, GND, MT11, T11_n, T12_n, T12, MT12, T12_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U2044(WL15_n, WL16, __A02_1__OVFSTB_n, WL15, WL16_n, __A02_3__UNF, GND,  ,  ,  ,  , __A02_3__OVF, __A02_1__OVFSTB_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U2045(__A02_3__OVF, OVF_n, __A02_3__UNF, UNF_n, __A02_2__SB0, __A02_2__SB0_n, GND, __A02_2__SB1_n, __A02_2__SB1, SB2_n, __A02_2__SB2, T12A, T12_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U2046(__A02_NET_158, P04, P05_n, __A02_NET_155, STOP_n, __A02_NET_156, GND, __A02_NET_157,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);


    U74HC02 #(1, 0, 0, 0) U3001(__A03_NET_166, NISQ, __A03_1__NISQL, __A03_NET_167, STRTFC, __A03_NET_168, GND, RT_n, __A03_NET_163, RBSQ, __A03_NET_163, WT_n, __A03_1__wsqg, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3002(__A03_NET_166, __A03_1__INKBT1, T12_n, __A03_NET_166, __A03_1__RPTFRC, __A03_NET_168, GND, __A03_1__CSQG, T12_n, CT_n, __A03_NET_167, __A03_1__NISQL, STRTFC, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(0, 1, 1, 0, 0, 1) U3003(__A03_1__NISQL, __A03_1__NISQL_n, __A03_NET_168, __A03_NET_163, __A03_1__wsqg, __A03_1__WSQG_n, GND, STRTFC, __A03_NET_161, __A03_1__SQEXT, __A03_NET_175, SQEXT_n, __A03_NET_174, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3004(__A03_NET_197, WL16_n, __A03_1__WSQG_n, __A03_NET_210, WL14_n, __A03_1__WSQG_n, GND, WL13_n, __A03_1__WSQG_n, __A03_NET_209,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U3005(__A03_NET_161, GOJAM, MTCSAI, __A03_NET_165, __A03_1__NISQL_n, T12_n, GND, STRTFC, __A03_NET_165, __A03_NET_172, __A03_NET_172, __A03_NET_164, __A03_NET_171, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U3006(EXTPLS, EXT, __A03_NET_164, __A03_1__INKBT1, STRTFC, FUTEXT, GND, __A03_NET_175, __A03_1__RPTFRC, __A03_NET_171, __A03_NET_174, __A03_NET_164, FUTEXT, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 1) U3007(__A03_NET_170, __A03_NET_172, FUTEXT, __A03_NET_174, __A03_NET_175, __A03_NET_170, GND, INHPLS, __A03_1__INHINT, __A03_NET_169, KRPT, __A03_1__IIP, __A03_1__IIP_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U3008(__A03_NET_175, __A03_1__MSQEXT, __A03_NET_169, __A03_1__MINHL, __A03_1__IIP_n, __A03_1__MIIP, GND, __A03_1__MSQ16, __A03_NET_202, __A03_1__MSQ14, __A03_NET_188, __A03_1__MSQ13, __A03_NET_190, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3009(__A03_NET_169, RELPLS, __A03_1__IIP_n, GOJAM, n5XP4, __A03_1__IIP, GND, __A03_NET_196, FUTEXT, __A03_1__NISQL_n, T12_n, __A03_1__INHINT, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3010(PHS2_n, RUPTOR_n, OVNHRP, __A03_1__INHINT, __A03_1__IIP, __A03_NET_194, GND, __A03_NET_192, __A03_NET_193, STRTFC, T02, __A03_NET_195, MNHRPT, VCC, SIM_RST, SIM_CLK);
    assign RPTSET = RPTSET_U3011_2;
    assign RPTSET = RPTSET_U3011_4;
    assign RPTSET = RPTSET_U3011_6;
    U74LVC07 U3011(__A03_NET_196, RPTSET_U3011_2, __A03_NET_195, RPTSET_U3011_4, __A03_NET_194, RPTSET_U3011_6, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 1, 1, 1) U3012(__A03_NET_193, RPTSET, __A03_NET_192, __A03_NET_202, __A03_NET_197, __A03_1__SQR16, GND, __A03_NET_210, __A03_1__SQR14, __A03_NET_188, __A03_NET_209, __A03_1__SQR13, __A03_NET_190, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3013(__A03_NET_202, __A03_1__RPTFRC, __A03_NET_188, __A03_1__RPTFRC, __A03_1__CSQG, __A03_1__SQR14, GND, __A03_1__SQR13, __A03_NET_190, __A03_1__RPTFRC, __A03_1__CSQG, __A03_1__SQR16, __A03_1__CSQG, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U3014(__A03_NET_200, __A03_NET_202, INKL, __A03_NET_199, INKL, __A03_1__SQR16, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U3015(__A03_NET_189, __A03_NET_187, __A03_NET_190, __A03_NET_187, __A03_NET_203, __A03_NET_201, GND, __A03_NET_208, __A03_NET_189, __A03_NET_188, __A03_NET_203, __A03_NET_198, __A03_NET_203, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3016(__A03_NET_190, __A03_NET_188, __A03_NET_189, __A03_NET_187, __A03_NET_186, __A03_NET_206, GND, __A03_NET_178, __A03_NET_190, __A03_NET_187, __A03_NET_186, __A03_NET_207, __A03_NET_203, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 0, 1) U3017(__A03_NET_189, __A03_NET_186, __A03_NET_190, __A03_NET_188, __A03_NET_186, __A03_NET_204, GND, __A03_NET_191, __A03_1__RPTFRC, __A03_NET_185, __A03_1__SQR12, __A03_NET_205, __A03_NET_188, VCC, SIM_RST, SIM_CLK);
    U74HC04 U3018(__A03_NET_201, SQ1_n, __A03_NET_208, SQ2_n, __A03_NET_207, __A03_1__SQ3_n, GND, __A03_1__SQ4_n, __A03_NET_206, __A03_1__SQ6_n, __A03_NET_205, __A03_1__SQ7_n, __A03_NET_204, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3019(__A03_NET_185, WL12_n, __A03_1__WSQG_n, __A03_NET_177, WL11_n, __A03_1__WSQG_n, GND, __A03_NET_191, __A03_1__CSQG, __A03_1__SQR12, __A03_NET_176, __A03_1__CSQG, __A03_1__SQR11, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 1, 0) U3020(__A03_1__RPTFRC, __A03_NET_177, __A03_1__RPTFRC, __A03_NET_184, __A03_NET_183, __A03_NET_182, GND, __A03_1__INKBT1, INKL, T01_n, STD2, __A03_NET_176, __A03_1__SQR11, VCC, SIM_RST, SIM_CLK);
    U74HC04 U3021(__A03_NET_191, __A03_1__MSQ12, __A03_NET_176, __A03_1__MSQ11, __A03_NET_182, __A03_1__MSQ10, GND, SQR12_n, __A03_1__SQR12, __A03_1__RPTFRC, __A03_NET_193, __A03_1__SQ5_n, __A03_NET_178, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3022(__A03_1__QC0, __A03_1__SQR11, __A03_1__SQR12, __A03_NET_181, __A03_NET_176, __A03_1__SQR12, GND, __A03_1__SQR11, __A03_NET_191, __A03_NET_180, __A03_NET_191, __A03_NET_176, __A03_NET_179, VCC, SIM_RST, SIM_CLK);
    U74HC04 U3023(__A03_1__QC0, QC0_n, __A03_NET_181, QC1_n, __A03_NET_180, QC2_n, GND, QC3_n, __A03_NET_179, SQR10, __A03_NET_182, SQR10_n, __A03_NET_183, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3024(__A03_NET_184, WL10_n, __A03_1__WSQG_n, __A03_NET_183, __A03_NET_182, __A03_1__CSQG, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U3025(__A03_NET_200, __A03_NET_186, __A03_NET_199, __A03_NET_203, __A03_NET_188, __A03_NET_187, GND, __A03_NET_189, __A03_NET_190, SQ0_n, __A03_NET_198, MP3A, MP3_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3026(__A03_NET_227, __A03_1__SQ5_n, QC0_n, __A03_NET_228, __A03_1__SQ5_n, SQEXT_n, GND, __A03_NET_227, __A03_NET_228, __A03_NET_229, __A03_NET_229, ST0_n, IC1, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(0, 0, 0, 0, 0, 1) U3027(__A03_NET_227, __A03_2__SQ5QC0_n, IC2, IC2_n, __A03_NET_233, EXST1_n, GND, TC0_n, TC0, IC3, __A03_2__IC3_n, __A03_2__NEXST0_n, __A03_2__NEXST0, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3028(IC2, __A03_NET_229, ST1_n, __A03_NET_226, SQEXT_n, __A03_1__QC0, GND, SQEXT_n, ST1_n, __A03_NET_233, __A03_NET_233, __A03_2__NEXST0, __A03_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3029(__A03_NET_226, __A03_1__SQ6_n, SQ1_n, __A03_2__NEXST0_n, __A03_1__QC0, TCF0, GND, __A03_2__IC3_n, TC0, STD2, TCF0, IC11, ST0_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3030(IC6, __A03_NET_232, __A03_1__SQ3_n, IC7, __A03_NET_232, __A03_1__SQ4_n, GND, SQ0_n, __A03_2__NEXST0_n, TC0, __A03_1__SQEXT, ST0_n, __A03_2__NEXST0, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3031(DCS0, __A03_1__SQ4_n, EXST0_n, DCA0, EXST0_n, __A03_1__SQ3_n, GND, DCS0, DCA0, __A03_2__IC4_n, QC1_n, ST1_n, __A03_NET_216, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3032(IC7, IC6, IC1, DCS0, DCA0, __A03_NET_220, GND, IC5, __A03_NET_214, __A03_1__SQ5_n, __A03_1__SQEXT, __A03_NET_221, IC11, VCC, SIM_RST, SIM_CLK);
    assign __A03_2__IC13_n = __A03_2__IC13_n_U3033_2;
    assign __A03_2__IC13_n = __A03_2__IC13_n_U3033_4;
    U74LVC07 U3033(__A03_NET_221, __A03_2__IC13_n_U3033_2, __A03_NET_220, __A03_2__IC13_n_U3033_4,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U3034(__A03_2__IC4_n, IC4, __A03_2__IC13_n, IC13, IC5, IC5_n, GND, IC9, __A03_2__IC9_n, QXCH0_n, __A03_2__QXCH0, EXST0_n, __A03_NET_213, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3035(__A03_NET_215, QC3_n, ST0_n, __A03_NET_214, __A03_NET_216, __A03_NET_215, GND, __A03_2__LXCH0, DXCH0, IC8_n, ST0_n, SQEXT_n, __A03_NET_213, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3036(__A03_2__NEXST0_n, QC1_n, SQ2_n, QC1_n, EXST0_n, __A03_2__QXCH0, GND, TS0, __A03_1__SQ5_n, QC2_n, __A03_2__NEXST0_n, __A03_2__LXCH0, SQ2_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U3037(__A03_2__IC9_n, IC5, TS0, __A03_2__QXCH0, __A03_2__LXCH0, __A03_NET_223, GND, __A03_NET_222, SQ2_n, QC0_n, __A03_1__SQEXT, ST1_n, __A03_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC04 U3038(TS0, TS0_n, IC10_n, IC10, DAS0, DAS0_n, GND, __A03_2__BZF0_n, __A03_2__BZF0, __A03_2__BMF0_n, __A03_2__BMF0, IC16, IC16_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3039(__A03_1__SQ5_n, __A03_2__NEXST0_n, SQ2_n, __A03_2__NEXST0_n, QC0_n, DAS0, GND, IC10_n, IC4, DXCH0, DAS0, DXCH0, QC1_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3040(SQ1_n, QC0_n, EXST0_n, QC0_n, __A03_1__SQ6_n, __A03_2__BMF0, GND, CCS0, SQ1_n, QC0_n, __A03_2__NEXST0_n, __A03_2__BZF0, EXST0_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3041(IC15_n, __A03_2__BMF0, __A03_2__BZF0, __A03_NET_218, __A03_2__BZF0_n, BR2_n, GND, __A03_2__BMF0_n, BR1B2B, __A03_NET_217, __A03_NET_218, __A03_NET_217, IC16_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U3042(IC17, IC16, IC15_n, DAS1_n, __A03_NET_212, ADS0, GND, CCS0, MSU0, IC12_n, __A03_1__SQ7_n, __A03_2__NEXST0_n, MASK0, VCC, SIM_RST, SIM_CLK);
    U74HC04 U3043(IC15_n, IC15, CCS0, CCS0_n, DAS1_n, DAS1, GND, IC12, IC12_n, MSU0_n, MSU0, AUG0_n, __A03_2__AUG0, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 0, 1) U3044(SQ2_n, QC3_n, QC2_n, SQ2_n, __A03_2__NEXST0_n, INCR0, GND, MSU0, SQ2_n, EXST0_n, QC0_n, ADS0, __A03_2__NEXST0_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3045(SQ2_n, EXST0_n, SQ2_n, EXST0_n, QC3_n, __A03_2__DIM0, GND, MP3, ST3_n, __A03_1__SQ7_n, SQEXT_n, __A03_2__AUG0, QC2_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(0, 0, 1, 0, 0, 0) U3046(__A03_2__DIM0, DIM0_n, MP3, MP3_n, MP1, MP1_n, GND, MP0_n, MP0, TCSAJ3_n, __A03_2__TCSAJ3, RSM3_n, RSM3, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3047(ST1_n, __A03_1__SQ7_n, ST0_n, __A03_1__SQ7_n, SQEXT_n, MP0, GND, __A03_2__TCSAJ3, SQ0_n, __A03_1__SQEXT, ST3_n, MP1, SQEXT_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3048(ST3_n, __A03_2__SQ5QC0_n, __A03_1__SQ6_n, EXST0_n, QC0_n, SU0, GND, __A03_NET_219, MP0, MASK0, RXOR0, RSM3, __A03_1__SQEXT, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(0, 0, 0, 0, 1, 0) U3049(MASK0, MASK0_n, __A03_NET_219, IC14, __A03_2__NDX0, NDX0_n, GND, NDXX1_n, __A03_2__NDXX1, GOJ1_n, GOJ1, IC11_n, IC11, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3050(AD0, __A03_2__NEXST0_n, __A03_1__SQ6_n,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U3051(__A03_2__NEXST0_n, __A03_1__SQ5_n, SQEXT_n, __A03_1__SQ5_n, ST1_n, __A03_2__NDXX1, GND, GOJ1, __A03_1__SQEXT, ST1_n, SQ0_n, __A03_2__NDX0, QC0_n, VCC, SIM_RST, SIM_CLK);


    U74HC02 #(0, 0, 0, 1) U4001(T12USE_n, DVST, __A04_NET_243, DIVSTG, T12USE_n, T03, GND, __A04_NET_244, __A04_NET_242, __A04_NET_268, GOJAM, MTCSAI, __A04_NET_249, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U4002(T03, T12USE_n, T12USE_n, RSTSTG, GOJAM, __A04_NET_243, GND, __A04_NET_242, PHS3_n, __A04_NET_243, T12_n, __A04_NET_244, PHS3_n, VCC, SIM_RST, SIM_CLK);
    assign __A04_NET_250 = __A04_NET_250_U4003_2;
    assign __A04_NET_250 = __A04_NET_250_U4003_4;
    assign __A04_NET_238 = __A04_NET_238_U4003_6;
    assign __A04_NET_238 = __A04_NET_238_U4003_8;
    assign __A04_1__SGUM = __A04_1__SGUM_U4003_10;
    assign __A04_1__SGUM = __A04_1__SGUM_U4003_12;
    U74LVC07 U4003(__A04_NET_249, __A04_NET_250_U4003_2, __A04_NET_248, __A04_NET_250_U4003_4, __A04_NET_229, __A04_NET_238_U4003_6, GND, __A04_NET_238_U4003_8, __A04_NET_232, __A04_1__SGUM_U4003_10, __A04_NET_198, __A04_1__SGUM_U4003_12, __A04_NET_197, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 1, 0) U4004(ST1, __A04_NET_245, __A04_1__STG1, __A04_1__STG3, __A04_1__STG2, __A04_NET_231, GND, __A04_NET_254, __A04_1__STG2, __A04_1__STG3, __A04_NET_236, __A04_NET_248, __A04_NET_247, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4005(__A04_NET_247, __A04_NET_250, T01, __A04_NET_245, __A04_NET_234, __A04_NET_269, GND, __A04_NET_268, __A04_NET_250, __A04_NET_241, __A04_NET_247, __A04_NET_268, __A04_NET_246, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U4006(__A04_NET_236, __A04_NET_241, __A04_1__STG1, __A04_1__STG1, __A04_NET_236, __A04_NET_246, GND, ST2, __A04_NET_230, __A04_NET_229, __A04_NET_234, __A04_NET_236, __A04_NET_235, VCC, SIM_RST, SIM_CLK);
    U74HC04 U4007(__A04_NET_236, __A04_1__MST1, __A04_NET_259, __A04_1__MST2, __A04_NET_269, __A04_1__MST3, GND, __A04_1__MBR1, __A04_NET_216, __A04_1__MBR2, __A04_NET_212, __A04_NET_234, DVST, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(0, 1, 1, 1, 0, 0) U4008(__A04_NET_231, ST0_n, __A04_NET_254, ST1_n, __A04_NET_264, ST3_n, GND, __A04_1__ST4_n, __A04_NET_252, __A04_1__ST376_n, __A04_1__ST376, DV1376_n, DV1376, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U4009(__A04_NET_235, MTCSAI, __A04_NET_238, GOJAM, T01, __A04_NET_233, GND, __A04_NET_264, __A04_1__STG3, __A04_NET_259, __A04_NET_236, __A04_NET_232, __A04_NET_233, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U4010(__A04_NET_230, __A04_NET_211, XT1_n, XB7_n, NDR100_n, __A04_NET_240, GND, __A04_NET_239, __A04_NET_256, STRTFC, T01, RSTSTG, __A04_NET_261, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U4011(__A04_NET_262, __A04_NET_268, __A04_NET_238, __A04_NET_237, __A04_NET_233, __A04_NET_268, GND, __A04_NET_262, __A04_1__STG2, __A04_NET_259, __A04_NET_259, __A04_NET_237, __A04_1__STG2, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U4012(__A04_NET_260, __A04_NET_234, __A04_NET_259, __A04_NET_256, __A04_NET_260, __A04_NET_261, GND, __A04_NET_268, __A04_NET_256, __A04_NET_265, __A04_NET_261, __A04_NET_268, __A04_NET_266, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 0, 0) U4013(__A04_NET_269, __A04_NET_265, __A04_1__STG3, __A04_1__STG3, __A04_NET_269, __A04_NET_266, GND, __A04_1__STG1, __A04_1__STG3, __A04_NET_251, __A04_NET_259, __A04_NET_251, __A04_1__ST376, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U4014(STD2, INKL, __A04_1__STG1, __A04_1__STG3, __A04_NET_259, __A04_NET_267, GND, __A04_NET_263, SQ0_n, EXST1_n, QC3_n, SQR10_n, RUPT1, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4015(__A04_NET_269, __A04_1__STG1, QC0_n, SQEXT_n, SQ1_n, __A04_NET_253, GND, __A04_NET_198, SUMB16_n, SUMA16_n, TSGU_n, __A04_NET_252, __A04_1__STG2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4016(__A04_NET_255, __A04_NET_252, __A04_1__ST376, __A04_1__DV3764, DIV_n, __A04_NET_255, GND, __A04_NET_254, __A04_1__ST376, __A04_1__ST1376_n, DIV_n, __A04_1__ST1376_n, DV1376, VCC, SIM_RST, SIM_CLK);
    U74HC04 U4017(__A04_NET_253, DIV_n, __A04_1__DV0, __A04_1__DV0_n, DV1, DV1_n, GND, DV376_n, __A04_1__DV376, __A04_NET_189, TL15, BR1, __A04_NET_216, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4018(__A04_1__DV0, DIV_n, ST0_n, DV1, DIV_n, ST1_n, GND, DIV_n, __A04_1__ST4_n, DV4, DIV_n, __A04_1__ST376_n, __A04_1__DV376, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4019(__A04_NET_183, SUMA16_n, SUMB16_n, __A04_NET_197, PHS4, PHS3_n, GND, UNF_n, TOV_n, __A04_NET_186, L15_n, __A04_NET_189, __A04_NET_191, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 0, 1) U4020(PHS4_n, WL16_n, __A04_NET_191, __A04_NET_188, __A04_NET_215, __A04_NET_194, GND, __A04_NET_195, __A04_NET_216, __A04_NET_193, __A04_NET_192, __A04_NET_188, TSGN_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4021(__A04_NET_193, TSGN_n, PHS3_n, __A04_NET_192, __A04_NET_189, PHS3_n, GND, TOV_n, PHS2_n, __A04_NET_205, __A04_1__SGUM, __A04_NET_186, __A04_NET_187, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U4022(__A04_NET_196, __A04_NET_183, PHS3_n, TSGU_n, PHS4, __A04_NET_184, GND, __A04_NET_185, WL16_n, WL15_n, WL14_n, WL13_n, __A04_NET_217, VCC, SIM_RST, SIM_CLK);
    assign __A04_NET_216 = __A04_NET_216_U4023_2;
    assign __A04_NET_216 = __A04_NET_216_U4023_4;
    assign __A04_NET_215 = __A04_NET_215_U4023_6;
    assign __A04_NET_215 = __A04_NET_215_U4023_8;
    assign __A04_NET_221 = __A04_NET_221_U4023_10;
    assign __A04_NET_221 = __A04_NET_221_U4023_12;
    U74LVC07 U4023(__A04_NET_187, __A04_NET_216_U4023_2, __A04_NET_194, __A04_NET_216_U4023_4, __A04_NET_195, __A04_NET_215_U4023_6, GND, __A04_NET_215_U4023_8, __A04_NET_190, __A04_NET_221_U4023_10, __A04_NET_217, __A04_NET_221_U4023_12, __A04_NET_220, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 0, 0) U4024(__A04_NET_190, __A04_NET_205, __A04_NET_196, __A04_NET_200, TOV_n, OVF_n, GND, __A04_NET_210, PHS3_n, __A04_NET_207, TMZ_n, PHS4_n, __A04_NET_222, VCC, SIM_RST, SIM_CLK);
    U74HC04 U4025(__A04_NET_215, BR1_n, __A04_1__TSGN2, __A04_NET_210, __A04_NET_212, BR2, GND, BR2_n, __A04_NET_204, DV4_n, DV4, __A04_NET_332, __A04_NET_331, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4026(GEQZRO_n, PHS4_n, WL16_n, PHS4_n, __A04_NET_210, __A04_NET_202, GND, __A04_NET_203, __A04_NET_202, __A04_NET_221, __A04_NET_204, __A04_NET_201, TPZG_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U4027(__A04_NET_220, WL12_n, WL11_n, WL10_n, WL09_n, __A04_NET_226, GND, __A04_NET_223, WL08_n, WL07_n, WL06_n, WL05_n, __A04_NET_219, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(0, 1) U4028(__A04_NET_218, WL04_n, WL03_n, WL02_n, WL01_n, __A04_NET_228, GND, __A04_NET_227, __A04_NET_212, __A04_NET_207, __A04_NET_206, __A04_NET_205, __A04_NET_204, VCC, SIM_RST, SIM_CLK);
    assign __A04_NET_221 = __A04_NET_221_U4029_2;
    assign __A04_NET_221 = __A04_NET_221_U4029_4;
    assign __A04_NET_221 = __A04_NET_221_U4029_6;
    assign __A04_NET_212 = __A04_NET_212_U4029_8;
    assign __A04_NET_212 = __A04_NET_212_U4029_10;
    U74LVC07 U4029(__A04_NET_219, __A04_NET_221_U4029_2, __A04_NET_218, __A04_NET_221_U4029_4, __A04_NET_222, __A04_NET_221_U4029_6, GND, __A04_NET_212_U4029_8, __A04_NET_199, __A04_NET_212_U4029_10, __A04_NET_203,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U4030(__A04_NET_206, TMZ_n, PHS3_n, __A04_NET_199, __A04_NET_201, __A04_NET_200, GND, SQ0_n, EXST0_n, __A04_NET_331, QC3_n, SQEXT_n, __A04_NET_277, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4031(__A04_NET_332, SQR10, QC0_n, __A04_NET_332, SQR10_n, __A04_2__WRITE0, GND, RAND0, SQR10, __A04_NET_332, QC1_n, READ0, QC0_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U4032(READ0, __A04_2__READ0_n, __A04_2__WRITE0, __A04_2__WRITE0_n, WOR0, __A04_2__WOR0_n, GND, RXOR0_n, RXOR0, __A04_2__RUPT0_n, RUPT0, __A04_2__RUPT1_n, RUPT1, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4033(QC1_n, SQR10_n, SQR10, __A04_NET_332, QC2_n, ROR0, GND, WOR0, QC2_n, __A04_NET_332, SQR10_n, WAND0, __A04_NET_332, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4034(SQR10, __A04_NET_332, QC3_n, __A04_NET_332, SQR10_n, RUPT0, GND, __A04_NET_275, ST0_n, SQR12_n, SQ2_n, RXOR0, QC3_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U4035(__A04_NET_275, __A04_NET_276, INOUT, INOUT_n, __A04_NET_280, __A04_NET_317, GND, BR1B2_n, __A04_2__BR1B2, BR12B_n, __A04_2__BR12B, BR1B2B_n, BR1B2B, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4036(PRINC, __A04_NET_277, __A04_NET_276, RRPA, T03_n, __A04_2__RUPT1_n, GND, T03_n, RXOR0_n, n3XP7, __A04_NET_270, T03_n, __A04_NET_273, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4037(EXST0_n, SQ0_n, INOUT, DV4, PRINC, __A04_NET_311, GND, __A04_NET_327, __A04_NET_273, __A04_NET_271, __A04_NET_278, INOUT, __A04_2__RUPT0_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4038(__A04_NET_270, ROR0, WOR0, __A04_NET_272, T03_n, __A04_NET_274, GND, RAND0, WAND0, __A04_NET_274, DV4_n, T05_n, n5XP28, VCC, SIM_RST, SIM_CLK);
    assign RB_n = RB_n_U4039_2;
    assign RC_n = RC_n_U4039_4;
    assign n5XP11 = n5XP11_U4039_6;
    assign n5XP11 = n5XP11_U4039_8;
    assign RA_n = RA_n_U4039_10;
    assign WG_n = WG_n_U4039_12;
    U74LVC07 U4039(__A04_NET_327, RB_n_U4039_2, __A04_NET_326, RC_n_U4039_4, __A04_NET_329, n5XP11_U4039_6, GND, n5XP11_U4039_8, __A04_NET_328, RA_n_U4039_10, __A04_NET_330, WG_n_U4039_12, __A04_NET_300, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4040(__A04_NET_272, __A04_NET_282, T05_n, INOUT_n, READ0, __A04_NET_329, GND, WCH_n, __A04_NET_283, n7XP14, __A04_NET_284, __A04_NET_326, __A04_NET_279, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4041(__A04_NET_328, __A04_2__WRITE0, RXOR0, __A04_NET_271, __A04_2__READ0_n, T05_n, GND, __A04_2__WRITE0_n, T05_n, __A04_NET_283, T05_n, __A04_2__WOR0_n, __A04_NET_284, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4042(__A04_NET_282, T05_n, RXOR0_n, __A04_NET_285, T02_n, __A04_2__WRITE0_n, GND, T02_n, INOUT_n, n2XP3, T09_n, __A04_2__RUPT0_n, n9XP1, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4043(__A04_NET_283, __A04_NET_282, RUPT1, IC13, IC12, __A04_NET_286, GND, __A04_NET_300, n9XP1, __A04_NET_279, __A04_NET_278, __A04_NET_330, n2XP3, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4044(__A04_NET_279, T09_n, RXOR0_n, __A04_NET_278, T09_n, __A04_NET_286, GND, __A04_NET_282, __A04_NET_285, __A04_NET_337, T01_n, __A04_2__RUPT1_n, RB2, VCC, SIM_RST, SIM_CLK);
    assign WG_n = WG_n_U4045_2;
    assign __A04_NET_280 = __A04_NET_280_U4045_4;
    assign __A04_NET_280 = __A04_NET_280_U4045_6;
    assign RA_n = RA_n_U4045_8;
    assign WG_n = WG_n_U4045_10;
    assign TMZ_n = TMZ_n_U4045_12;
    U74LVC07 U4045(__A04_NET_337, WG_n_U4045_2, __A04_NET_335, __A04_NET_280_U4045_4, __A04_NET_336, __A04_NET_280_U4045_6, GND, RA_n_U4045_8, __A04_NET_314, WG_n_U4045_10, __A04_NET_301, TMZ_n_U4045_12, __A04_NET_323, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4046(RUPT0, RUPT1, INOUT, MP1, MP3A, __A04_NET_335, GND, __A04_NET_336, __A04_1__DV0, IC15, DV1376, __A04_NET_281, RSM3, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4047(R15, __A04_NET_281, T01_n, n1XP10, T01_n, __A04_1__DV0_n, GND, MP0_n, T03_n, __A04_NET_288, INOUT_n, T03_n, __A04_NET_319, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4048(T02_n, __A04_1__DV0_n, BRDIF_n, TS0_n, T04_n, __A04_NET_299, GND, __A04_NET_294, T04_n, BR1, MP0_n, n2XP5, BR1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4049(n3XP2, T03_n, TS0_n, __A04_2__BR1B2, BR1, BR2_n, GND, BR1_n, BR2, __A04_2__BR12B, __A04_2__BR1B2, __A04_2__BR12B, BRDIF_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4050(BR1B2B, BR2, BR1, n4XP5, TS0_n, T04_n, GND, T04_n, INOUT_n, n4XP11, T04_n, MP3_n, __A04_NET_324, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4051(MP0_n, BR1_n, DV1_n, T04_n, BR2_n, __A04_NET_289, GND, __A04_NET_293, TS0_n, T05_n, BR1B2_n, __A04_NET_321, T04_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4052(T05_n, TS0_n, T07_n, BR1_n, MP3_n, n7XP19, GND, n8XP6, T08_n, DV1_n, BR2, __A04_NET_309, BR12B_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4053(B15X, T05_n, DV1_n, n5XP4, T05_n, RSM3_n, GND, T06_n, DV1_n, n6XP5, T06_n, MP3_n, TL15, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4054(__A04_1__TSGN2, T07_n, MP0_n, __A04_NET_308, T07_n, DV1_n, GND, T08_n, DV1_n, n8XP5, T09_n, MP3_n, __A04_NET_313, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4055(T09_n, BR1, T09_n, MP0_n, BR1_n, __A04_NET_296, GND, __A04_NET_298, MP0_n, T09_n, BRDIF_n, __A04_NET_318, MP0_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4056(KRPT, T09_n, __A04_2__RUPT1_n, MP0T10, T10_n, MP0_n, GND, __A04_NET_317, T02_n, __A04_NET_315, STORE1_n, T09_n, __A04_NET_303, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4057(MP3_n, MP0_n, n1XP10, n8XP5, __A04_NET_313, __A04_NET_314, GND,  ,  ,  ,  , __A04_NET_316, T11_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U4058(RSC_n, __A04_2__MRSC, __A04_NET_316, __A04_NET_312, TRSM, __A04_NET_211, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 1) U4059( ,  , __A04_NET_319, B15X, n7XP19, __A04_NET_325, GND, __A04_NET_320, n8XP5, __A04_NET_318, __A04_NET_296,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U4060(__A04_NET_323, n2XP5, n1XP10, __A04_NET_291, __A04_NET_299, __A04_NET_298, GND, n1XP10, MP0T10, __A04_NET_290, __A04_NET_293, __A04_NET_316, __A04_NET_292, VCC, SIM_RST, SIM_CLK);
    assign WY_n = WY_n_U4061_2;
    assign WY_n = WY_n_U4061_4;
    assign WL_n = WL_n_U4061_6;
    assign RC_n = RC_n_U4061_8;
    assign RB_n = RB_n_U4061_10;
    assign CI_n = CI_n_U4061_12;
    U74LVC07 U4061(__A04_NET_325, WY_n_U4061_2, __A04_NET_320, WY_n_U4061_4, __A04_NET_322, WL_n_U4061_6, GND, RC_n_U4061_8, __A04_NET_297, RB_n_U4061_10, __A04_NET_295, CI_n_U4061_12, __A04_NET_291, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U4062(__A04_NET_294, __A04_NET_321, __A04_NET_321, n2XP5, __A04_NET_296, __A04_NET_297, GND, __A04_NET_295, __A04_NET_294, n7XP19, __A04_NET_318, __A04_NET_322, n6XP5, VCC, SIM_RST, SIM_CLK);
    assign TSGN_n = TSGN_n_U4063_2;
    assign TSGN_n = TSGN_n_U4063_4;
    assign RB1_n = RB1_n_U4063_6;
    assign __A04_2__L16_n = __A04_2__L16_n_U4063_8;
    assign R1C_n = R1C_n_U4063_10;
    assign n8PP4 = n8PP4_U4063_12;
    U74LVC07 U4063(__A04_NET_290, TSGN_n_U4063_2, __A04_NET_287, TSGN_n_U4063_4, __A04_NET_292, RB1_n_U4063_6, GND, __A04_2__L16_n_U4063_8, __A04_NET_312, R1C_n_U4063_10, __A04_NET_310, n8PP4_U4063_12, __A04_NET_311, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4064(__A04_NET_289, __A04_NET_288,  ,  ,  ,  , GND,  ,  ,  ,  , __A04_NET_287, __A04_NET_308, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4065(__A04_NET_310, __A04_NET_316, __A04_NET_309, __A04_2__BRXP3, T03_n, IC15_n, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC4002 U4066(RSC_n, __A04_NET_315, __A04_NET_324, __A04_NET_308, __A04_2__BRXP3, __A04_NET_307, GND, __A04_NET_306, __A04_NET_315, __A04_NET_303, __A04_NET_324, __A04_2__BRXP3, __A04_NET_301, VCC, SIM_RST, SIM_CLK);


    U74HC27 U5001(IC10, IC3, TC0, TCF0, IC4, __A05_NET_249, GND, __A05_NET_248, IC2, IC3, RSM3, __A05_NET_251, IC2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5002(__A05_NET_250, STD2, IC2, __A05_NET_270, T01_n, __A05_NET_251, GND, T01_n, __A05_NET_250, __A05_NET_253, IC10_n, T01_n, __A05_NET_247, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5003(__A05_NET_266, T01_n, __A05_NET_249, __A05_NET_252, T02_n, __A05_NET_248, GND, T08_n, CCS0_n, __A05_NET_206, T02_n, MP3_n, n2XP7, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U5004(T02_n, STD2, __A05_1__10XP6, __A05_1__10XP7, __A05_NET_247, __A05_NET_256, GND, __A05_NET_259, __A05_NET_253, n3XP6, __A05_NET_243, DVST, DIV_n, VCC, SIM_RST, SIM_CLK);
    assign MONEX_n = MONEX_n_U5005_2;
    assign RZ_n = RZ_n_U5005_4;
    assign RB_n = RB_n_U5005_6;
    assign RA_n = RA_n_U5005_8;
    assign WA_n = WA_n_U5005_10;
    assign RL_n = RL_n_U5005_12;
    U74LVC07 U5005(__A05_NET_256, MONEX_n_U5005_2, __A05_NET_259, RZ_n_U5005_4, __A05_NET_260, RB_n_U5005_6, GND, RA_n_U5005_8, __A05_NET_258, WA_n_U5005_10, __A05_NET_246, RL_n_U5005_12, __A05_NET_240, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5006(__A05_NET_252, __A05_1__8XP15, __A05_NET_242, __A05_NET_241, __A05_1__8XP12, __A05_NET_240, GND, __A05_1__PARTC, INKL_n, SHIFT, MONPCH, __A05_1__NISQ_n, n2XP7, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5007(__A05_1__3XP5, T03_n, IC2_n, __A05_NET_274, T01_n, IC15_n, GND, __A05_NET_274, __A05_NET_276, __A05_NET_258, T03_n, TC0_n, n3XP6, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5008(__A05_NET_276, T04_n, IC2_n, __A05_NET_244, T02_n, IC15_n, GND, __A05_NET_244, __A05_NET_275, TPZG_n, T04_n, DAS0_n, __A05_NET_242, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 0, 0) U5009(__A05_NET_246, __A05_NET_242, __A05_NET_245, __A05_NET_245, T04_n, MASK0_n, GND, MP3_n, T10_n, __A05_NET_241, T05_n, IC2_n, __A05_NET_243, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5010(__A05_NET_275, T05_n, __A05_NET_255, __A05_NET_254, __A05_NET_274, __A05_NET_275, GND, T05_n, DAS0_n, n5XP12, T06_n, RSM3_n, __A05_NET_279, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5011(__A05_1__PARTC, PRINC, __A05_NET_275, __A05_NET_274, n7XP9, __A05_NET_227, GND, __A05_NET_278, n9XP5, __A05_NET_274, __A05_NET_279, __A05_NET_255, CCS0, VCC, SIM_RST, SIM_CLK);
    assign TMZ_n = TMZ_n_U5012_2;
    assign WG_n = WG_n_U5012_4;
    assign RG_n = RG_n_U5012_6;
    assign RC_n = RC_n_U5012_8;
    assign A2X_n = A2X_n_U5012_10;
    assign WY_n = WY_n_U5012_12;
    U74LVC07 U5012(__A05_NET_254, TMZ_n_U5012_2, __A05_NET_278, WG_n_U5012_4, __A05_NET_281, RG_n_U5012_6, GND, RC_n_U5012_8, __A05_NET_277, A2X_n_U5012_10, __A05_NET_262, WY_n_U5012_12, __A05_NET_264, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5013(__A05_NET_280, T06_n, DAS0_n, __A05_NET_263, T06_n, MSU0_n, GND, __A05_NET_245, __A05_NET_263, __A05_NET_277, T07_n, DAS0_n, __A05_NET_265, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 1) U5014(__A05_NET_275, __A05_NET_261, __A05_NET_261, __A05_NET_280, __A05_NET_263, __A05_NET_262, GND, __A05_NET_264, __A05_NET_261, __A05_NET_263, __A05_NET_280, __A05_NET_281, __A05_NET_280, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U5015(__A05_NET_260, __A05_NET_266, __A05_1__3XP5, __A05_NET_265, __A05_NET_279, __A05_NET_268, GND, __A05_NET_267, IC3, RSM3, MP3, IC16, TSUDO_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5016(n7XP9, T07_n, MSU0_n, __A05_NET_261, T07_n, IC2_n, GND, T07_n, CCS0_n, __A05_NET_271, __A05_NET_203, __A05_NET_195, __A05_NET_202, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 0, 1) U5017(__A05_NET_263, __A05_NET_270, __A05_1__8XP3, __A05_NET_271, n4XP5, __A05_NET_273, GND, __A05_NET_269, n4XP5, __A05_NET_271, __A05_NET_270, __A05_NET_272, __A05_1__10XP6, VCC, SIM_RST, SIM_CLK);
    assign CI_n = CI_n_U5018_2;
    assign RZ_n = RZ_n_U5018_4;
    assign WY12_n = WY12_n_U5018_6;
    assign WZ_n = WZ_n_U5018_8;
    assign RB_n = RB_n_U5018_10;
    assign WB_n = WB_n_U5018_12;
    U74LVC07 U5018(__A05_NET_272, CI_n_U5018_2, __A05_NET_273, RZ_n_U5018_4, __A05_NET_269, WY12_n_U5018_6, GND, WZ_n_U5018_8, __A05_NET_205, RB_n_U5018_10, __A05_NET_202, WB_n_U5018_12, __A05_NET_213, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 0, 1) U5019(CCS0_n, T07_n, BR1_n, CCS0_n, T07_n, PTWOX, GND, __A05_NET_205, __A05_1__3XP5, __A05_NET_192, __A05_NET_206, n7XP4, BR2_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5020(INKL_n, FETCH0, __A05_NET_206, __A05_NET_208, n9XP5, __A05_NET_210, GND, __A05_NET_207, IC2, IC4, DXCH0, __A05_NET_203, T08_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U5021(RAD, TSUDO_n, T08_n, __A05_NET_213, RAD, __A05_NET_197, GND, T08_n, __A05_NET_212, __A05_1__8XP15, T08_n, __A05_NET_209, __A05_1__8XP3, VCC, SIM_RST, SIM_CLK);
    U74HC04 U5022(IC16, __A05_NET_212, __A05_NET_289, RQ_n, MP3, __A05_NET_299, GND, SCAD_n, SCAD, NDR100_n, __A05_NET_292, __A05_NET_336, __A05_NET_329, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5023(__A05_NET_209, MP0, IC1, __A05_NET_208, T08_n, __A05_NET_207, GND, T08_n, __A05_NET_196, __A05_NET_197, T08_n, GOJ1_n, __A05_1__RSTRT, VCC, SIM_RST, SIM_CLK);
    assign RU_n = RU_n_U5024_2;
    assign RA_n = RA_n_U5024_4;
    assign ST2_n = ST2_n_U5024_6;
    assign WY_n = WY_n_U5024_8;
    assign RC_n = RC_n_U5024_10;
    assign WA_n = WA_n_U5024_12;
    U74LVC07 U5024(__A05_NET_210, RU_n_U5024_2, __A05_NET_200, RA_n_U5024_4, __A05_NET_198, ST2_n_U5024_6, GND, WY_n_U5024_8, __A05_NET_235, RC_n_U5024_10, __A05_NET_237, WA_n_U5024_12, __A05_NET_219, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5025(DXCH0, GOJ1, T08_n, BR2, T10_n, __A05_1__10XP6, GND, __A05_NET_199, IC1, IC10, RUPT0, __A05_NET_196, DAS0, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5026(__A05_1__8XP12, T08_n, DAS0_n, __A05_NET_192, T08_n, TCSAJ3_n, GND, T09_n, __A05_NET_194, __A05_NET_195, IC2, __A05_1__DV1B1B, __A05_NET_194, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5027(n9XP5, T09_n, DAS0_n, __A05_NET_230, T09_n, MASK0_n, GND, __A05_NET_230, __A05_NET_234, __A05_NET_200, T10_n, T08_n, __A05_NET_231, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5028(__A05_NET_198, __A05_NET_192, __A05_NET_231, n10XP1, __A05_NET_199, T10_n, GND, T10_n, __A05_NET_229, __A05_NET_234, DAS0, __A05_NET_239, __A05_NET_229, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U5029(__A05_NET_231, __A05_NET_230, T10_n, DAS0_n, BR1B2_n, n10XP8, GND, __A05_NET_219, __A05_NET_195, __A05_NET_220, n5XP11, __A05_NET_235, __A05_NET_234, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5030(__A05_NET_239, MSU0_n, BR1_n, __A05_1__10XP7, T10_n, __A05_NET_232, GND, __A05_NET_239, __A05_NET_233, __A05_NET_232, BR12B_n, DAS0_n, __A05_NET_233, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5031(n11XP2, T11_n, MSU0_n, __A05_NET_236, T10_n, MASK0_n, GND, __A05_NET_230, __A05_NET_236, __A05_NET_237, T10_n, __A05_NET_238, __A05_NET_220, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5032(__A05_NET_238, MSU0, IC14, __A05_NET_221, INCSET_n, __A05_NET_217, GND, GOJAM, __A05_1__GHNHC, __A05_NET_228, __A05_NET_228, T01, __A05_1__GHNHC, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U5033(__A05_NET_218, C24A, C25A, C26A, C27A, __A05_NET_225, GND, __A05_NET_224, C30A, C37P, C40P, C41P, __A05_NET_216, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 0, 1) U5034(C42P, C43P, IC12, DAS0, DAS1, __A05_NET_355, GND, __A05_NET_351, RL10BB, __A05_NET_310, __A05_2__RSCT, __A05_NET_215, C44P, VCC, SIM_RST, SIM_CLK);
    assign __A05_NET_217 = __A05_NET_217_U5035_2;
    assign __A05_NET_217 = __A05_NET_217_U5035_4;
    assign __A05_NET_217 = __A05_NET_217_U5035_6;
    assign __A05_NET_311 = __A05_NET_311_U5035_8;
    assign __A05_NET_311 = __A05_NET_311_U5035_10;
    assign WS_n = WS_n_U5035_12;
    U74LVC07 U5035(__A05_NET_218, __A05_NET_217_U5035_2, __A05_NET_216, __A05_NET_217_U5035_4, __A05_NET_215, __A05_NET_217_U5035_6, GND, __A05_NET_311_U5035_8, __A05_NET_355, __A05_NET_311_U5035_10, __A05_NET_354, WS_n_U5035_12, __A05_NET_351, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5036(__A05_1__PINC_n, __A05_NET_221, PINC, PINC, __A05_1__PINC_n, T12, GND, T01_n, __A05_NET_311, RL10BB, T01_n, FETCH0_n, R6, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U5037(__A05_NET_354, IC9, DXCH0, PRINC, INOUT, __A05_NET_353, GND, __A05_NET_352, YB0_n, YT0_n, S12, S11, __A05_NET_292, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5038(__A05_NET_310, T01_n, CHINC_n, __A05_NET_286, T03_n, __A05_NET_313, GND, IC5, MP0, __A05_NET_356, T03_n, IC8_n, __A05_NET_312, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 0, 1) U5039(T01_n, MONPCH, TS0, DAS0, MASK0, __A05_NET_359, GND, __A05_NET_357, __A05_NET_286, __A05_NET_312, __A05_NET_289, __A05_2__RSCT, INKL_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U5040(__A05_NET_287, __A05_NET_290,  ,  ,  ,  , GND,  ,  ,  ,  , __A05_NET_358, __A05_2__6XP2, VCC, SIM_RST, SIM_CLK);
    assign WB_n = WB_n_U5041_2;
    assign WB_n = WB_n_U5041_4;
    assign __A05_NET_313 = __A05_NET_313_U5041_6;
    assign __A05_NET_313 = __A05_NET_313_U5041_8;
    assign RL_n = RL_n_U5041_10;
    assign RA_n = RA_n_U5041_12;
    U74LVC07 U5041(__A05_NET_357, WB_n_U5041_2, __A05_NET_358, WB_n_U5041_4, __A05_NET_359, __A05_NET_313_U5041_6, GND, __A05_NET_313_U5041_8, __A05_NET_356, RL_n_U5041_10, __A05_NET_346, RA_n_U5041_12, __A05_NET_347, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5042(n2XP8, T02_n, FETCH0_n, __A05_NET_289, T03_n, QXCH0_n, GND, T04_n, DV1_n, __A05_NET_288, T04_n, __A05_NET_291, __A05_NET_287, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5043(__A05_NET_312, __A05_NET_288, DV1, INOUT, IC2, __A05_NET_291, GND, __A05_NET_345, __A05_NET_290, __A05_NET_285, __A05_2__5XP9, __A05_NET_346, __A05_2__11XP6, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5044(__A05_NET_347, __A05_NET_286, __A05_2__6XP2, TRSM, T05_n, NDX0_n, GND, IC12_n, T05_n, __A05_NET_290, DAS1_n, T05_n, __A05_NET_285, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 0, 1) U5045(__A05_2__5XP13, n5XP15, DAS1, PRINC, __A05_1__PARTC, __A05_NET_282, GND, __A05_NET_350, __A05_NET_283, n2XP8, __A05_2__10XP10, __A05_NET_344, __A05_NET_297, VCC, SIM_RST, SIM_CLK);
    assign RG_n = RG_n_U5046_2;
    assign RG_n = RG_n_U5046_4;
    assign WY_n = WY_n_U5046_6;
    assign A2X_n = A2X_n_U5046_8;
    assign CI_n = CI_n_U5046_10;
    assign WY12_n = WY12_n_U5046_12;
    U74LVC07 U5046(__A05_NET_345, RG_n_U5046_2, __A05_NET_344, RG_n_U5046_4, __A05_NET_350, WY_n_U5046_6, GND, A2X_n_U5046_8, __A05_NET_348, CI_n_U5046_10, __A05_NET_349, WY12_n_U5046_12, __A05_NET_372, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U5047(__A05_NET_283, __A05_NET_282, T05_n, __A05_NET_348, __A05_NET_285, __A05_2__10XP10, GND, SHIFT_n, T05_n, __A05_2__5XP9, SHANC_n, T05_n, __A05_NET_284, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5048(__A05_NET_284, __A05_NET_298, YT0_n, YB0_n, XT0_n, __A05_NET_373, GND, __A05_NET_296, RAND0, WAND0, __A05_NET_329, __A05_NET_349, __A05_NET_300, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5049(__A05_2__5XP13, IC8_n, T05_n, n5XP15, QXCH0_n, T05_n, GND, CHINC_n, T05_n, n5XP21, IC5_n, T05_n, __A05_NET_297, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U5050(__A05_NET_298, IC16_n, T05_n, __A05_NET_300, __A05_NET_299, T05_n, GND, __A05_NET_298, __A05_NET_300, __A05_NET_372, S11, S12, __A05_NET_374, VCC, SIM_RST, SIM_CLK);
    assign RB_n = RB_n_U5051_2;
    assign RZ_n = RZ_n_U5051_4;
    assign SCAD = SCAD_U5051_6;
    assign SCAD = SCAD_U5051_8;
    assign RC_n = RC_n_U5051_10;
    assign __A05_NET_330 = __A05_NET_330_U5051_12;
    U74LVC07 U5051(__A05_NET_371, RB_n_U5051_2, __A05_NET_370, RZ_n_U5051_4, __A05_NET_374, SCAD_U5051_6, GND, SCAD_U5051_8, __A05_NET_373, RC_n_U5051_10, __A05_NET_363, __A05_NET_330_U5051_12, __A05_NET_361, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5052(__A05_NET_371, __A05_2__5XP19, __A05_NET_298, __A05_NET_370, __A05_2__6XP7, __A05_NET_300, GND, XT2_n, NDR100_n, OCTAD2, NDR100_n, XT3_n, __A05_2__OCTAD3, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5053(__A05_2__OCTAD4, NDR100_n, XT4_n, __A05_2__OCTAD5, NDR100_n, XT5_n, GND, NDR100_n, XT6_n, __A05_2__OCTAD6, BR1_n, DV1_n, __A05_NET_329, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5054(__A05_NET_295, __A05_NET_296, T05_n, __A05_2__5XP19, T05_n, __A05_NET_294, GND, DV1_n, BR1, __A05_1__DV1B1B, TS0_n, BRDIF_n, __A05_NET_331, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(0, 1) U5055(__A05_NET_363, __A05_NET_295, __A05_NET_333, __A05_NET_324, __A05_NET_323, __A05_NET_362, GND, __A05_NET_364, __A05_2__5XP13, __A05_NET_308, __A05_NET_340, __A05_NET_317, __A05_NET_338, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5056(ROR0, __A05_1__DV1B1B, IC2, IC5, READ0, __A05_NET_361, GND, __A05_NET_365, IC2, IC3, TS0, __A05_NET_294, WOR0, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 0, 1) U5057(__A05_NET_360, __A05_NET_331, DV4, __A05_NET_334, __A05_NET_330, T05_n, GND, __A05_NET_336, T05_n, __A05_NET_335, __A05_NET_334, __A05_NET_333, __A05_NET_368, VCC, SIM_RST, SIM_CLK);
    assign __A05_NET_330 = __A05_NET_330_U5058_2;
    assign __A05_2__Z16_n = __A05_2__Z16_n_U5058_4;
    assign WA_n = WA_n_U5058_6;
    assign __A05_NET_332 = __A05_NET_332_U5058_8;
    assign __A05_NET_332 = __A05_NET_332_U5058_10;
    assign WZ_n = WZ_n_U5058_12;
    U74LVC07 U5058(__A05_NET_360, __A05_NET_330_U5058_2, __A05_NET_369, __A05_2__Z16_n_U5058_4, __A05_NET_368, WA_n_U5058_6, GND, __A05_NET_332_U5058_8, __A05_NET_365, __A05_NET_332_U5058_10, __A05_NET_366, WZ_n_U5058_12, __A05_NET_367, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(0, 1, 0, 0, 0, 0) U5059(__A05_NET_335, __A05_NET_369, __A05_NET_328, __A05_NET_367, __A05_NET_333, __A05_NET_343, GND, __A05_NET_322, __A05_NET_324, NISQ, __A05_1__NISQ_n, __A05_1__MNISQ, __A05_1__NISQ_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5060(__A05_NET_366, IC16, MP3, __A05_NET_328, T06_n, __A05_NET_332, GND, T06_n, DAS1_n, n6XP8, n6XP8, __A05_2__6XP7, __A05_NET_306, VCC, SIM_RST, SIM_CLK);
    assign TOV_n = TOV_n_U5061_2;
    assign RU_n = RU_n_U5061_4;
    assign RU_n = RU_n_U5061_6;
    assign WB_n = WB_n_U5061_8;
    assign RG_n = RG_n_U5061_10;
    assign TSGN_n = TSGN_n_U5061_12;
    U74LVC07 U5061(__A05_NET_306, TOV_n_U5061_2, __A05_NET_303, RU_n_U5061_4, __A05_NET_302, RU_n_U5061_6, GND, WB_n_U5061_8, __A05_NET_304, RG_n_U5061_10, __A05_NET_314, TSGN_n_U5061_12, __A05_NET_342, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5062(__A05_2__6XP7, DV4_n, T06_n, __A05_NET_316, T07_n, __A05_NET_305, GND, T07_n, STFET1_n, __A05_NET_315, T08_n, DV4_n, RSTSTG, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5063(__A05_NET_328, n6XP8, __A05_NET_309, __A05_NET_340, __A05_NET_308, __A05_NET_302, GND, __A05_2__6XP2, T06_n, RXOR0, INOUT_n, __A05_NET_303, n5XP11, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U5064(IC13, IC14, __A05_NET_316, __A05_NET_340, __A05_NET_309, __A05_NET_304, GND, __A05_NET_314, __A05_NET_316, __A05_NET_315, __A05_NET_323, __A05_NET_305, DV1, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5065(T08_n, MONWBK, IC2, IC14, DV1, __A05_NET_321, GND, __A05_NET_318, DV4B1B, IC4, __A05_NET_320, U2BBK, STFET1_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5066(__A05_NET_342, RSTSTG, __A05_2__5XP9, __A05_NET_333, T09_n, __A05_NET_336, GND, T09_n, DV4_n, __A05_NET_340, T09_n, DAS1_n, __A05_NET_324, VCC, SIM_RST, SIM_CLK);
    assign __A05_2__Z15_n = __A05_2__Z15_n_U5067_2;
    assign WL_n = WL_n_U5067_4;
    assign TMZ_n = TMZ_n_U5067_6;
    assign WYD_n = WYD_n_U5067_8;
    assign TSGN_n = TSGN_n_U5067_10;
    U74LVC07 U5067(__A05_NET_343, __A05_2__Z15_n_U5067_2, __A05_NET_338, WL_n_U5067_4, __A05_NET_322, TMZ_n_U5067_6, GND, WYD_n_U5067_8, __A05_NET_326, TSGN_n_U5067_10, __A05_NET_227,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U5068(__A05_NET_309, T10_n, __A05_NET_321,  ,  ,  , GND, T10_n, IC11_n, __A05_2__10XP10, T10_n, __A05_NET_318, __A05_NET_317, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5069(DAS1_n, ADS0, T12_n, T12USE_n, DV1_n, __A05_NET_308, GND,  ,  ,  ,  , __A05_NET_320, BR2, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U5070(DV4B1B, DV4_n, BR1, __A05_2__11XP6, T11_n, DV1_n, GND, __A05_2__5XP9, __A05_2__11XP6, __A05_NET_326, T11_n, RXOR0_n, __A05_NET_323, VCC, SIM_RST, SIM_CLK);


    U74HC27 U6001(T04, T07, __A06_NET_284, __A06_NET_285, __A06_NET_286, __A06_NET_283, GND, __A06_NET_301, T01, T03, T05, __A06_NET_298, T10, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6002(__A06_NET_284, __A06_NET_298, DV376_n, __A06_NET_285, T01_n, DV1376_n, GND, T04_n, DV4_n, __A06_NET_286, MP1_n, __A06_NET_287, __A06_NET_288, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 0, 1) U6003(T07, T09, __A06_1__L15A_n, __A06_1__L02A_n, L01_n, __A06_NET_300, GND, __A06_NET_341, T05, T08, T11, __A06_NET_302, T11, VCC, SIM_RST, SIM_CLK);
    assign __A06_NET_287 = __A06_NET_287_U6004_2;
    assign __A06_NET_287 = __A06_NET_287_U6004_4;
    assign A2X_n = A2X_n_U6004_6;
    assign RB_n = RB_n_U6004_8;
    assign WYD_n = WYD_n_U6004_10;
    assign WY_n = WY_n_U6004_12;
    U74LVC07 U6004(__A06_NET_301, __A06_NET_287_U6004_2, __A06_NET_302, __A06_NET_287_U6004_4, __A06_NET_299, A2X_n_U6004_6, GND, RB_n_U6004_8, __A06_NET_313, WYD_n_U6004_10, __A06_NET_314, WY_n_U6004_12, __A06_NET_305, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 1, 1, 0) U6005(__A06_NET_312, __A06_NET_288, n2XP7, L2GD_n, __A06_1__ZIP, __A06_1__DVXP1, GND, __A06_1__DVXP1, __A06_NET_306, __A06_NET_314, __A06_NET_303, __A06_NET_304, __A06_NET_307, VCC, SIM_RST, SIM_CLK);
    U74HC04 U6006(L01_n, __A06_NET_290, __A06_1__L02A_n, __A06_NET_340, __A06_1__L15A_n, __A06_NET_289, GND, __A06_1__DVXP1, __A06_NET_283, __A06_1__ZIP, __A06_NET_312, __A06_NET_338, __A06_NET_339, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U6007(n7XP19, __A06_1__ZIP, __A06_1__DVXP1, __A06_NET_309, RBSQ, __A06_NET_313, GND, __A06_NET_316, __A06_NET_290, __A06_NET_340, __A06_NET_289, __A06_NET_299, __A06_1__DVXP1, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6008(__A06_NET_289, __A06_NET_290, __A06_NET_312, __A06_NET_304, __A06_NET_303, __A06_NET_315, GND, __A06_NET_339, __A06_NET_303, __A06_NET_304, __A06_1__L02A_n, __A06_NET_304, __A06_1__L02A_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6009(__A06_NET_306, __A06_NET_312, __A06_NET_307, __A06_NET_311, __A06_NET_312, __A06_NET_338, GND, __A06_NET_341, DV376_n, __A06_NET_310, DV1376_n, T02_n, __A06_NET_272, VCC, SIM_RST, SIM_CLK);
    U74HC04 U6010(__A06_NET_311, MCRO_n, __A06_NET_277, __A06_NET_274, __A06_NET_281, __A06_NET_282, GND, __A06_1__ZAP, ZAP_n, __A06_NET_343, __A06_NET_341, MONEX, MONEX_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6011(__A06_NET_312, __A06_NET_338, __A06_NET_339, __A06_NET_316, __A06_NET_312, __A06_NET_309, GND, __A06_NET_303, __A06_NET_340, __A06_1__L15A_n, L01_n, __A06_1__ZIPCI, __A06_NET_300, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 1, 1, 0) U6012(__A06_NET_277, __A06_NET_310, __A06_NET_272, __A06_NET_281, __A06_NET_276, DIVSTG, GND, T08, T10, __A06_NET_278, MP1_n, __A06_NET_280, __A06_NET_266, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U6013(T06, T09, DV376_n, __A06_NET_275, T12USE_n, __A06_NET_276, GND, __A06_NET_279, T02, T04, T06, __A06_NET_275, T12, VCC, SIM_RST, SIM_CLK);
    assign __A06_NET_280 = __A06_NET_280_U6014_2;
    assign __A06_NET_280 = __A06_NET_280_U6014_4;
    assign WL_n = WL_n_U6014_6;
    assign RG_n = RG_n_U6014_8;
    assign WB_n = WB_n_U6014_10;
    assign RU_n = RU_n_U6014_12;
    U74LVC07 U6014(__A06_NET_279, __A06_NET_280_U6014_2, __A06_NET_278, __A06_NET_280_U6014_4, __A06_NET_273, WL_n_U6014_6, GND, RG_n_U6014_8, __A06_NET_270, WB_n_U6014_10, __A06_NET_291, RU_n_U6014_12, __A06_NET_292, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 1, 0) U6015(__A06_NET_268, T01, T03, __A06_NET_267, __A06_NET_268, MP3_n, GND, __A06_NET_266, __A06_NET_267, ZAP_n, n5XP28, __A06_NET_274, TSGU_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 1, 1, 0) U6016(__A06_NET_273, __A06_NET_274, n5XP12, __A06_NET_297, RRPA, n5XP4, GND, n5XP15, n3XP6, WQ_n, n9XP5, n6XP8, __A06_NET_346, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(0, 1) U6017(__A06_NET_270, n5XP4, RADRG, __A06_NET_274, n5XP28, __A06_NET_271, GND, __A06_NET_269, n5XP28, n1XP10, __A06_NET_282, n2XP3, __A06_NET_291, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U6018(__A06_NET_292, __A06_NET_282, __A06_1__ZAP, n5XP12, n6XP5, __A06_NET_293, GND, __A06_NET_294, PRINC, PINC, MINC, DINC, __A06_NET_229, VCC, SIM_RST, SIM_CLK);
    assign WZ_n = WZ_n_U6019_2;
    assign TOV_n = TOV_n_U6019_4;
    assign WSC_n = WSC_n_U6019_6;
    assign WG_n = WG_n_U6019_8;
    assign __A06_NET_217 = __A06_NET_217_U6019_10;
    assign __A06_NET_217 = __A06_NET_217_U6019_12;
    U74LVC07 U6019(__A06_NET_297, WZ_n_U6019_2, __A06_NET_345, TOV_n_U6019_4, __A06_NET_346, WSC_n_U6019_6, GND, WG_n_U6019_8, __A06_NET_342, __A06_NET_217_U6019_10, __A06_NET_218, __A06_NET_217_U6019_12, __A06_NET_219, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6020(n6XP5, n3XP2, BR1_n, PHS4_n, TSGU_n, __A06_1__RB1F, GND, CLXC, TSGU_n, BR1, PHS4_n, __A06_NET_345, n9XP5, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 1, 1) U6021(__A06_NET_342, n6XP8, n6XP8, PIFL_n, __A06_1__DVXP1, __A06_NET_344, GND, PTWOX, MONEX, __A06_NET_327, MONEX, B15X, __A06_NET_328, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6022(PIFL_n, __A06_NET_343, STBE, n1XP10, STBF, __A06_NET_326, GND, __A06_NET_218, __A06_NET_263, __A06_NET_262, INCR0, __A06_NET_344, T02, VCC, SIM_RST, SIM_CLK);
    U74HC04 U6023(__A06_NET_327, TWOX, __A06_NET_328, BXVX, __A06_NET_336, __A06_NET_317, GND, __A06_NET_319, __A06_NET_317, __A06_NET_325, __A06_NET_319, __A06_NET_324, __A06_NET_325, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6024(CGMC, __A06_NET_326, __A06_NET_336, __A06_NET_318, CGMC, __A06_NET_321, GND, __A06_NET_318, __A06_NET_326, __A06_NET_336, BR1, AUG0_n, __A06_NET_263, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(0, 0, 0, 0, 1, 0) U6025(__A06_NET_324, __A06_NET_323, __A06_NET_323, __A06_NET_320, __A06_NET_320, __A06_NET_322, GND, __A06_NET_321, __A06_NET_322, __A06_NET_210, __A06_NET_212, __A06_NET_225, __A06_2__7XP10, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6026(__A06_NET_262, DIM0_n, BR12B_n, __A06_NET_219, PINC, __A06_NET_261, GND, BR12B_n, DINC_n, __A06_NET_261, T06_n, __A06_NET_217, __A06_2__6XP10, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6027(__A06_NET_222, MINC, MCDU, __A06_NET_220, AUG0_n, BR1_n, GND, DIM0_n, BR1B2B_n, __A06_NET_221, BR1B2B_n, DINC_n, __A06_NET_211, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6028(__A06_NET_220, __A06_NET_221, BR1B2B_n, CDUSTB_n, DINC_n, __A06_2__POUT, GND, __A06_2__MOUT, BR12B_n, CDUSTB_n, DINC_n, __A06_NET_216, __A06_NET_211, VCC, SIM_RST, SIM_CLK);
    assign __A06_NET_223 = __A06_NET_223_U6029_2;
    assign __A06_NET_223 = __A06_NET_223_U6029_4;
    assign MONEX_n = MONEX_n_U6029_6;
    assign WA_n = WA_n_U6029_8;
    assign RB1_n = RB1_n_U6029_10;
    assign R1C_n = R1C_n_U6029_12;
    U74LVC07 U6029(__A06_NET_222, __A06_NET_223_U6029_2, __A06_NET_216, __A06_NET_223_U6029_4, __A06_NET_210, MONEX_n_U6029_6, GND, WA_n_U6029_8, __A06_NET_234, RB1_n_U6029_10, __A06_NET_225, R1C_n_U6029_12, __A06_NET_224, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6030(__A06_NET_212, T06_n, __A06_NET_223, __A06_NET_213, PCDU, MCDU, GND, T06_n, __A06_NET_213, __A06_2__6XP12, __A06_NET_233, T07_n, __A06_NET_235, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 1) U6031(BR2_n, DINC_n, DAS0, DAS1, MSU0, __A06_NET_233, GND, __A06_NET_234, __A06_NET_235, __A06_2__7XP7, __A06_NET_207, __A06_2__ZOUT, CDUSTB_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6032(__A06_NET_232, DV4_n, BR1B2B, __A06_2__7XP7, T07_n, __A06_NET_237, GND, WAND0, INOTLD, __A06_NET_240, T07_n, __A06_NET_240, n7XP14, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6033(__A06_NET_232, WAND0, DAS1_n, T07_n, BR1B2_n, __A06_2__7XP10, GND, __A06_2__7XP11, DAS1_n, T07_n, BR12B_n, __A06_NET_237, RAND0, VCC, SIM_RST, SIM_CLK);
    U74HC04 U6034(__A06_2__7XP11, __A06_NET_224, __A06_NET_201, PONEX, ST2_n, ST2, GND, ST1, __A06_NET_253, __A06_NET_250, __A06_2__PSEUDO, __A06_NET_251, __A06_2__RDBANK, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6035(__A06_2__7XP15, __A06_NET_230, T07_n, __A06_NET_239, __A06_NET_229, T07_n, GND, PRINC, INKL, __A06_NET_186, IC9, DXCH0, __A06_NET_187, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6036(PCDU, MCDU, n7XP9, n11XP2, __A06_2__7XP15, RUS_n, GND, __A06_NET_188, __A06_NET_239, __A06_NET_241, __A06_NET_207, __A06_NET_230, SHIFT, VCC, SIM_RST, SIM_CLK);
    assign RU_n = RU_n_U6037_2;
    assign WSC_n = WSC_n_U6037_4;
    assign WG_n = WG_n_U6037_6;
    assign RB_n = RB_n_U6037_8;
    assign n8PP4 = n8PP4_U6037_10;
    assign n8PP4 = n8PP4_U6037_12;
    U74LVC07 U6037(__A06_NET_188, RU_n_U6037_2, __A06_NET_189, WSC_n_U6037_4, __A06_NET_190, WG_n_U6037_6, GND, RB_n_U6037_8, __A06_NET_182, n8PP4_U6037_10, __A06_NET_181, n8PP4_U6037_12, __A06_NET_185, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6038(__A06_NET_186, T07_n, T04_n, MON_n, FETCH1, __A06_NET_191, GND, __A06_NET_189, __A06_2__WOVR, __A06_NET_191, __A06_NET_192, __A06_2__WOVR, MONPCH, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6039(__A06_NET_190, __A06_2__WOVR, __A06_NET_192, __A06_NET_192, T07_n, __A06_NET_187, GND, __A06_2__10XP9, __A06_NET_192, __A06_NET_182, T08_n, n8PP4, __A06_2__8XP4, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6040(RUPT1, DAS1, IC17, MASK0, IC11, __A06_NET_185, GND, __A06_NET_184, IC6, IC7, IC9, __A06_NET_181, MSU0, VCC, SIM_RST, SIM_CLK);
    assign n8PP4 = n8PP4_U6041_2;
    assign __A06_NET_203 = __A06_NET_203_U6041_4;
    assign __A06_NET_203 = __A06_NET_203_U6041_6;
    assign WS_n = WS_n_U6041_8;
    assign __A06_NET_206 = __A06_NET_206_U6041_10;
    assign __A06_NET_206 = __A06_NET_206_U6041_12;
    U74LVC07 U6041(__A06_NET_184, n8PP4_U6041_2, __A06_NET_204, __A06_NET_203_U6041_4, __A06_NET_202, __A06_NET_203_U6041_6, GND, WS_n_U6041_8, __A06_NET_205, __A06_NET_206_U6041_10, __A06_NET_195, __A06_NET_206_U6041_12, __A06_NET_194, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U6042(T08_n, RUPT0, __A06_NET_203, R6, R15, __A06_NET_205, GND, __A06_NET_194, ADS0, IC11, __A06_NET_193, __A06_NET_204, DAS0, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6043(__A06_NET_202, MP1, DV1376, __A06_NET_209, MP3_n, BR1_n, GND, __A06_NET_209, CCS0, __A06_NET_195, T11_n, __A06_NET_206, __A06_NET_207, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6044(__A06_NET_193, DAS1_n, BR2_n, __A06_NET_196, __A06_1__ZIPCI, __A06_2__6XP12, GND, CCS0_n, BR1B2B_n, __A06_NET_245, T10_n, NDXX1_n, EXT, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U6045(T03_n, DAS1_n, __A06_NET_248, __A06_NET_241, n2XP5, __A06_NET_260, GND, __A06_NET_257, IC7, DCS0, SU0, __A06_NET_241, ADS0, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1, 0) U6046(__A06_NET_201, n8XP6, n7XP4, n10XP8, __A06_2__6XP10, __A06_NET_199, GND, __A06_NET_200, IC6, DCA0, AD0, __A06_NET_245, __A06_NET_246, VCC, SIM_RST, SIM_CLK);
    assign CI_n = CI_n_U6047_2;
    assign WA_n = WA_n_U6047_4;
    assign RC_n = RC_n_U6047_6;
    assign __A06_NET_243 = __A06_NET_243_U6047_8;
    assign __A06_NET_243 = __A06_NET_243_U6047_10;
    assign ST2_n = ST2_n_U6047_12;
    U74LVC07 U6047(__A06_NET_196, CI_n_U6047_2, __A06_NET_260, WA_n_U6047_4, __A06_NET_258, RC_n_U6047_6, GND, __A06_NET_243_U6047_8, __A06_NET_257, __A06_NET_243_U6047_10, __A06_NET_256, ST2_n_U6047_12, __A06_NET_259, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6048(__A06_2__10XP9, T10_n, __A06_NET_246, __A06_NET_247, IC6, IC7, GND, T10_n, __A06_NET_247, __A06_NET_248, T10_n, __A06_NET_243, __A06_NET_242, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6049(__A06_NET_258, __A06_NET_242, __A06_2__7XP7, __A06_NET_256, __A06_NET_244, DV4B1B, GND, CCS0_n, BR12B_n, __A06_NET_244, T10_n, MP1_n, __A06_2__10XP15, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6050(__A06_2__8XP4, __A06_2__10XP15, __A06_2__8XP4, RADRZ, n9XP1, __A06_NET_252, GND, NEAC, __A06_NET_254, TL15, GOJAM, __A06_NET_259, RADRZ, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U6051(__A06_NET_253, n2XP8, n10XP1, MP0T10, __A06_2__10XP15, __A06_NET_334, GND, __A06_NET_264, __A06_1__DVXP1, GOJAM, NISQ, __A06_1__WHOMP_n, WHOMP, VCC, SIM_RST, SIM_CLK);
    assign RZ_n = RZ_n_U6052_2;
    assign RPTSET = RPTSET_U6052_4;
    assign RU_n = RU_n_U6052_6;
    assign RC_n = RC_n_U6052_8;
    U74LVC07 U6052(__A06_NET_252, RZ_n_U6052_2, __A06_NET_250, RPTSET_U6052_4, __A06_NET_251, RU_n_U6052_6, GND, RC_n_U6052_8, __A06_NET_335,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 0, 0) U6053(__A06_NET_254, MP0T10, NEAC, __A06_NET_249, RADRZ, __A06_2__PSEUDO, GND, T06_n, STFET1_n, __A06_2__RDBANK, __A06_1__ZIPCI, n3XP7, __A06_NET_335, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U6054(__A06_NET_249, GOJAM, n3XP7, n5XP21, n4XP11, RCH_n, GND,  ,  ,  ,  , __A06_2__PSEUDO, RADRG, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(0, 0, 0, 1, 0, 0) U6055(R1C_n, R1C, RB1_n, RB1, L02_n, __A06_NET_330, GND, __A06_1__L02A_n, __A06_NET_330, __A06_NET_329, L15_n, __A06_1__L15A_n, __A06_NET_329, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1, 0, 0, 0, 0, 0) U6056(__A06_NET_315, __A06_NET_305, __A06_1__WHOMP_n, WHOMPA,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 0, 0) U6057(__A06_1__WHOMP_n, WHOMP, CLXC,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);


    U74HC02 #(0, 1, 0, 0) U7001(__A07_1__WALSG, ZAP_n, WT_n, __A07_NET_166, __A07_NET_165, __A07_NET_167, GND, __A07_NET_166, WT_n, __A07_NET_169, WY_n, WT_n, __A07_NET_168, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1, 0, 0, 1, 1, 0) U7002(__A07_1__WALSG, WALSG_n, WY12_n, __A07_NET_165, WY_n, __A07_NET_167, GND, WYLOG_n, __A07_NET_169, WYHIG_n, __A07_NET_168, __A07_1__MWYG, __A07_NET_160, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 0, 1) U7003(__A07_NET_160, __A07_NET_169, __A07_NET_158, __A07_NET_158, WYD_n, WT_n, GND, __A07_NET_160, CT_n, CUG, L15_n, PIFL_n, __A07_NET_164, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1, 1, 1, 0, 0, 1) U7004(__A07_NET_158, WYDG_n, __A07_NET_162, WYDLOG_n, __A07_NET_163, WBG_n, GND, __A07_1__MWBG, WBG_n, __A07_1__MWG, __A07_1__WGA_n, WG1G_n, __A07_1__WGNORM, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 0, 1) U7005(__A07_NET_159, WYD_n, WT_n, __A07_NET_163, WB_n, WT_n, GND, WBG_n, CT_n, CBG, __A07_1__WGNORM, __A07_NET_175, WG2G_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U7006(SHIFT, NEAC, __A07_1__WGA_n, WT_n, GINH, __A07_1__WGNORM, GND, __A07_NET_175, __A07_1__WGA_n, WT_n, SR_n, __A07_NET_161, __A07_NET_164, VCC, SIM_RST, SIM_CLK);
    assign __A07_NET_162 = __A07_NET_162_U7007_2;
    assign __A07_NET_162 = __A07_NET_162_U7007_4;
    U74LVC07 U7007(__A07_NET_159, __A07_NET_162_U7007_2, __A07_NET_161, __A07_NET_162_U7007_4,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U7008(__A07_1__WGA_n, WT_n, __A07_1__WGA_n, WT_n, CYL_n, __A07_NET_170, GND, __A07_NET_174, __A07_1__WGA_n, WT_n, EDOP_n, __A07_NET_171, CYR_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U7009(__A07_NET_171, WG5G_n, __A07_NET_170, WG3G_n, __A07_NET_174, WEDOPG_n, GND, __A07_1__MWZG, WZG_n, __A07_1__MWLG, WLG_n, __A07_1__MWAG, WAG_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 0, 1) U7010(WG4G_n, __A07_NET_175, __A07_NET_171, __A07_NET_172, WT_n, WZ_n, GND, __A07_1__WSCG_n, XB5_n, __A07_NET_173, __A07_NET_172, __A07_NET_173, WZG_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7011(CZG, WZG_n, CT_n, __A07_NET_142, WL_n, WT_n, GND, __A07_1__WSCG_n, XB1_n, __A07_NET_145, __A07_NET_138, CT_n, CLG1G, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U7012(XB1_n, XT0_n, __A07_NET_142, __A07_NET_148, __A07_NET_145, WLG_n, GND, __A07_NET_139, __A07_NET_140, __A07_NET_141, __A07_1__WALSG, __A07_NET_148, __A07_1__WCHG_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U7013(__A07_NET_137, __A07_NET_142, __A07_NET_148, __A07_NET_145, __A07_1__WALSG, __A07_NET_143, GND, __A07_NET_144, __A07_NET_145, __A07_NET_148, __A07_NET_142, __A07_2__G2LSG, __A07_NET_138, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 0, 1) U7014(CLG2G, __A07_NET_137, CT_n, __A07_NET_140, WT_n, WA_n, GND, __A07_1__WSCG_n, XB0_n, __A07_NET_141, __A07_NET_140, __A07_NET_141, WAG_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7015(CAG, __A07_NET_139, CT_n, __A07_NET_155, WT_n, WS_n, GND, WSG_n, CT_n, CSG, WT_n, WQ_n, __A07_NET_154, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1, 0, 0, 0, 0, 1) U7016(__A07_NET_155, WSG_n, WSG_n, __A07_1__MWSG, WQG_n, __A07_1__MWQG, GND, __A07_1__P04A, P04_n, RCG_n, __A07_NET_209, G2LSG_n, __A07_2__G2LSG, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U7017(__A07_NET_154, __A07_NET_157, XB2_n, XT0_n, __A07_1__WCHG_n, __A07_NET_156, GND, __A07_1__PIPSAM_n, PIPPLS_n, SB2_n, __A07_1__P04A, WQG_n, __A07_NET_156, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7018(__A07_NET_157, __A07_1__WSCG_n, XB2_n, CQG, WQG_n, CT_n, GND, RT_n, RC_n, __A07_NET_209, RT_n, RQ_n, __A07_NET_210, VCC, SIM_RST, SIM_CLK);
    U74HC27 U7019(__A07_NET_210, __A07_NET_207, XB2_n, XT0_n, __A07_2__RCHG_n, __A07_NET_208, GND, __A07_2__RFBG_n, __A07_NET_213, __A07_NET_214, __A07_2__RBBK, RQG_n, __A07_NET_208, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7020(__A07_NET_207, __A07_2__RSCG_n, XB2_n, __A07_NET_213, __A07_2__RSCG_n, XB4_n, GND, __A07_2__RSCG_n, XB6_n, __A07_NET_214, __A07_NET_214, __A07_2__RBBK, __A07_2__RBBEG_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7021(__A07_2__G2LSG, TT_n, ZAP_n, __A07_NET_211, TT_n, L2GD_n, GND, TT_n, A2X_n, __A07_NET_205, T10_n, STFET1_n, __A07_2__RBBK, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1, 1, 0, 0, 0, 0) U7022(__A07_NET_211, L2GDG_n, __A07_NET_205, A2XG_n, __A07_NET_183, CGG, GND, __A07_2__MWEBG, __A07_2__WEBG_n, __A07_2__MWFBG, __A07_2__WFBG_n, __A07_2__WBBEG_n, __A07_NET_189, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7023(__A07_NET_204, L2GD_n, CT_n, __A07_NET_206, CT_n, WG_n, GND, __A07_1__WSCG_n, XB3_n, __A07_2__WEBG_n, __A07_NET_184, CT_n, __A07_2__CEBG, VCC, SIM_RST, SIM_CLK);
    U74HC27 U7024(__A07_NET_204, __A07_NET_206, __A07_2__WEBG_n, U2BBK, __A07_NET_189, __A07_NET_184, GND, __A07_NET_185, __A07_NET_189, U2BBK, __A07_NET_182, __A07_NET_183, CGMC, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7025(__A07_2__CFBG, __A07_NET_185, CT_n, __A07_NET_182, __A07_1__WSCG_n, T10_n, GND, __A07_NET_182, __A07_NET_189, __A07_2__WFBG_n, __A07_1__WSCG_n, XB6_n, __A07_NET_189, VCC, SIM_RST, SIM_CLK);
    U74HC04 U7026(__A07_2__WBBEG_n, __A07_2__MWBBEG, __A07_NET_190, RGG_n, RGG_n, __A07_2__MRGG, GND, __A07_2__MRAG, RAG_n, __A07_2__MRLG, RLG_n, __A07_2__REBG_n, __A07_NET_181, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7027(__A07_NET_190, RT_n, RG_n, __A07_NET_191, RT_n, RA_n, GND, __A07_NET_191, __A07_NET_186, RAG_n, XB0_n, __A07_2__RSCG_n, __A07_NET_186, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7028(__A07_NET_187, RT_n, RL_n, __A07_NET_188, __A07_2__RSCG_n, XB1_n, GND, RT_n, RZ_n, __A07_NET_178, __A07_NET_178, __A07_NET_177, RZG_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U7029(__A07_NET_187, __A07_NET_188, XB1_n, XT0_n, __A07_2__RCHG_n, __A07_NET_179, GND, US2SG, __A07_2__RUSG_n, SUMA15_n, SUMB15_n, RLG_n, __A07_NET_179, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7030(__A07_NET_177, XB5_n, __A07_2__RSCG_n, __A07_NET_181, __A07_2__RSCG_n, XB3_n, GND, RT_n, RU_n, __A07_NET_198, RT_n, RUS_n, __A07_NET_180, VCC, SIM_RST, SIM_CLK);
    U74HC04 U7031(__A07_NET_198, RUG_n, __A07_NET_180, __A07_2__RUSG_n, RULOG_n, __A07_2__MRULOG, GND, RBHG_n, __A07_NET_203, __A07_NET_201, RL10BB,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U7032(RULOG_n, __A07_NET_198, __A07_NET_180, __A07_NET_203, RT_n, RB_n, GND, RT_n, __A07_NET_201, __A07_NET_202, __A07_NET_203, __A07_NET_202, RBLG_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U7037( ,  ,  ,  ,  ,  , GND, __A07_NET_200, CI_n, __A07_1__WSCG_n, __A07_NET_149, __A07_2__RSCG_n, __A07_NET_196, VCC, SIM_RST, SIM_CLK);
    U74HC27 U7038( ,  , NEAC, EAC_n, MP3A, __A07_2__CINORM, GND, __A07_NET_196, RT_n, RSC_n, SCAD_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U7039(__A07_NET_199, __A07_NET_200, __A07_2__CIFF, __A07_2__CIFF, __A07_NET_199, CUG, GND, __A07_2__CIFF, __A07_2__CINORM, CI01_n, WSC_n, SCAD_n, __A07_NET_149, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7040(__A07_NET_197, RT_n, RCH_n, __A07_NET_153, WT_n, WCH_n, GND, WCH_n, CT_n, __A07_NET_151,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 #(0, 0, 0, 0, 1, 0) U7041(__A07_NET_197, __A07_2__RCHG_n, __A07_NET_153, __A07_1__WCHG_n, __A07_NET_151, __A07_1__CCHG_n, GND, __A07_NET_152, WG_n, __A07_1__WGA_n, __A07_NET_152, __A07_2__U2BBKG_n, U2BBK, VCC, SIM_RST, SIM_CLK);


    U74HC02 U8001(__A08_NET_205, A2XG_n, __A08_1___A1_n, __A08_NET_200, WYLOG_n, WL01_n, GND, WL16_n, WYDLOG_n, __A08_NET_199, __A08_1__Y1_n, CUG, __A08_1__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U8002(PONEX, __A08_NET_205, __A08_1__X1_n, CLXC, CUG, __A08_1__X1, GND, __A08_1__Y1_n, __A08_NET_200, __A08_NET_199, __A08_1__Y1, __A08_1__X1_n, __A08_1__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8003(__A08_NET_209, __A08_1__X1_n, __A08_1__Y1_n, XUY01_n, __A08_1__X1, __A08_1__Y1, GND, __A08_NET_209, XUY01_n, __A08_NET_207, __A08_NET_209, __A08_1___SUMA1, __A08_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8004( ,  , __A08_1___SUMA1, __A08_1___SUMB1, RULOG_n, __A08_NET_187, GND, __A08_NET_191, __A08_2___XUY1, XUY01_n, CI01_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U8005(CI01_n, __A08_NET_206, G01_n, __A08_1___GEM1, __A08_1___RL1_n, __A08_1___WL1, GND, WL01_n, __A08_1___WL1, __A08_1___MWL1, __A08_1___RL1_n, __A08_NET_157, __A08_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8006(__A08_1___SUMB1, __A08_NET_207, __A08_NET_206, __A08_NET_190, WAG_n, WL01_n, GND, WL03_n, WALSG_n, __A08_NET_192, __A08_1___A1_n, CAG, __A08_NET_188, VCC, SIM_RST, SIM_CLK);
    assign __A08_2___CO_IN = __A08_2___CO_IN_U8007_2;
    assign __A08_1___RL1_n = __A08_1___RL1_n_U8007_4;
    assign L01_n = L01_n_U8007_6;
    assign __A08_1___Z1_n = __A08_1___Z1_n_U8007_8;
    assign __A08_1___RL1_n = __A08_1___RL1_n_U8007_10;
    assign __A08_1___RL1_n = __A08_1___RL1_n_U8007_12;
    U74LVC07 U8007(__A08_NET_191, __A08_2___CO_IN_U8007_2, __A08_NET_185, __A08_1___RL1_n_U8007_4, __A08_NET_198, L01_n_U8007_6, GND, __A08_1___Z1_n_U8007_8, __A08_NET_221, __A08_1___RL1_n_U8007_10, __A08_NET_222, __A08_1___RL1_n_U8007_12, __A08_NET_220, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8008(__A08_NET_186, RAG_n, __A08_1___A1_n, __A08_NET_189, WLG_n, WL01_n, GND, __A08_2___G2_n, G2LSG_n, __A08_NET_196, L01_n, CLG1G, __A08_NET_197, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U8009( ,  ,  , __A08_NET_194, WQG_n, WL01_n, GND, __A08_NET_194, __A08_NET_193, __A08_1___Q1_n, __A08_1___Q1_n, CQG, __A08_NET_193, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U8010(__A08_NET_195, RQG_n, __A08_1___Q1_n, __A08_NET_224, WZG_n, WL01_n, GND, __A08_NET_224, __A08_NET_223, __A08_NET_221, __A08_1___Z1_n, CZG, __A08_NET_223, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8011(__A08_1___RL_OUT_1, __A08_NET_195, MDT01, RB1, R15, __A08_NET_220, GND, __A08_NET_227, __A08_NET_225, __A08_NET_226, __A08_NET_212, __A08_NET_222, __A08_NET_219, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U8012(__A08_NET_219, RZG_n, __A08_1___Z1_n, __A08_NET_228, WBG_n, WL01_n, GND, __A08_NET_228, __A08_NET_229, __A08_1___B1_n, __A08_1___B1_n, CBG, __A08_NET_229, VCC, SIM_RST, SIM_CLK);
    assign __A08_2___CO_IN = __A08_2___CO_IN_U8013_2;
    assign __A08_1___RL1_n = __A08_1___RL1_n_U8013_4;
    assign G01_n = G01_n_U8013_6;
    assign G01_n = G01_n_U8013_8;
    assign __A08_1___RL2_n = __A08_1___RL2_n_U8013_10;
    assign L02_n = L02_n_U8013_12;
    U74LVC07 U8013(__A08_NET_170, __A08_2___CO_IN_U8013_2, __A08_NET_227, __A08_1___RL1_n_U8013_4, __A08_NET_211, G01_n_U8013_6, GND, G01_n_U8013_8, __A08_NET_210, __A08_1___RL2_n_U8013_10, __A08_NET_137, L02_n_U8013_12, __A08_NET_147, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8014(__A08_NET_225, RBLG_n, __A08_1___B1_n, __A08_NET_226, __A08_NET_229, RCG_n, GND, WL16_n, WG3G_n, __A08_NET_216, WL02_n, WG4G_n, __A08_NET_215, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U8015(__A08_NET_190, __A08_NET_192, __A08_NET_187, __A08_NET_186, CH01, __A08_NET_185, GND, __A08_NET_198, __A08_NET_189, __A08_NET_196, __A08_NET_197, __A08_1___A1_n, __A08_NET_188, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8016(__A08_NET_214, L2GDG_n, MCRO_n, __A08_NET_213, WG1G_n, WL01_n, GND, G01_n, CGG, G01, RGG_n, G01_n, __A08_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U8017(__A08_NET_214, __A08_NET_213, WHOMPA, __A08_2___XUY2, XUY02_n, __A08_NET_170, GND, __A08_1___RL_OUT_1, RLG_n, L01_n, GND, __A08_NET_210, G01, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1, 0) U8018(__A08_NET_211, G01ED, SA01, __A08_NET_216, __A08_NET_215, __A08_NET_218, GND, __A08_NET_217, G02ED, SA02, __A08_NET_164, __A08_NET_163, __A08_NET_162, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8019(__A08_NET_158, A2XG_n, __A08_1___A2_n, __A08_NET_160, WYLOG_n, WL02_n, GND, WL01_n, WYDG_n, __A08_NET_159, __A08_1__Y2_n, CUG, __A08_1__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U8020(TWOX, __A08_NET_158, __A08_1__X2_n, CLXC, CUG, __A08_1__X2, GND, __A08_1__Y2_n, __A08_NET_160, __A08_NET_159, __A08_1__Y2, __A08_1__X2_n, __A08_1__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8021(__A08_NET_152, __A08_1__X2_n, __A08_1__Y2_n, XUY02_n, __A08_1__X2, __A08_1__Y2, GND,  ,  ,  , __A08_NET_152, XUY02_n, __A08_NET_155, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8022( ,  , __A08_NET_152, __A08_1___SUMA2, GND, __A08_2___CI_IN, GND, __A08_NET_156, __A08_1___SUMA2, __A08_1___SUMB2, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U8023(__A08_1___SUMB2, __A08_NET_155, __A08_NET_157, __A08_NET_141, WAG_n, WL02_n, GND, WL04_n, WALSG_n, __A08_NET_140, __A08_1___A2_n, CAG, __A08_NET_139, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U8024(__A08_NET_141, __A08_NET_140, __A08_NET_156, __A08_NET_142, CH02, __A08_NET_137, GND, __A08_NET_147, __A08_NET_175, __A08_NET_176, __A08_NET_177, __A08_1___A2_n, __A08_NET_139, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8025(__A08_NET_142, RAG_n, __A08_1___A2_n, __A08_NET_175, WLG_n, WL02_n, GND, G05_n, G2LSG_n, __A08_NET_176, L02_n, CLG1G, __A08_NET_177, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8026(RLG_n, L02_n, __A08_1___RL_OUT_2, __A08_NET_143, __A08_NET_149, __A08_NET_148, GND, __A08_NET_138, MDT02, R1C, RB2, __A08_1___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U8027(__A08_NET_179, WQG_n, WL02_n, __A08_1___Q2_n, __A08_NET_179, __A08_NET_178, GND, __A08_1___Q2_n, CQG, __A08_NET_178, RQG_n, __A08_1___Q2_n, __A08_NET_143, VCC, SIM_RST, SIM_CLK);
    assign __A08_1___RL2_n = __A08_1___RL2_n_U8028_2;
    assign __A08_1___Z2_n = __A08_1___Z2_n_U8028_4;
    assign __A08_1___RL2_n = __A08_1___RL2_n_U8028_6;
    assign __A08_1___RL2_n = __A08_1___RL2_n_U8028_8;
    assign __A08_1___G2_n = __A08_1___G2_n_U8028_10;
    assign __A08_1___G2_n = __A08_1___G2_n_U8028_12;
    U74LVC07 U8028(__A08_NET_148, __A08_1___RL2_n_U8028_2, __A08_NET_145, __A08_1___Z2_n_U8028_4, __A08_NET_138, __A08_1___RL2_n_U8028_6, GND, __A08_1___RL2_n_U8028_8, __A08_NET_180, __A08_1___G2_n_U8028_10, __A08_NET_162, __A08_1___G2_n_U8028_12, __A08_NET_169, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U8029(__A08_NET_144, WZG_n, WL02_n, __A08_NET_145, __A08_NET_144, __A08_NET_146, GND, __A08_1___Z2_n, CZG, __A08_NET_146, RZG_n, __A08_1___Z2_n, __A08_NET_149, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U8030(__A08_NET_183, WBG_n, WL02_n, __A08_1___B2_n, __A08_NET_183, __A08_NET_184, GND, __A08_1___B2_n, CBG, __A08_NET_184, RBLG_n, __A08_1___B2_n, __A08_NET_182, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U8031(__A08_NET_182, __A08_NET_181, __A08_NET_168, __A08_NET_167, G02, __A08_NET_169, GND, __A08_NET_263, GND, XUY06_n, __A08_2___XUY2, __A08_NET_180, __A08_NET_161, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8032(__A08_NET_181, __A08_NET_184, RCG_n, __A08_NET_164, WL01_n, WG3G_n, GND, WL03_n, WG4G_n, __A08_NET_163, L2GDG_n, L01_n, __A08_NET_168, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8033(__A08_NET_167, WG1G_n, WL02_n, G02, __A08_1___G2_n, CGG, GND, RGG_n, __A08_1___G2_n, __A08_NET_161,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U8034(__A08_1___G2_n, __A08_1___GEM2, __A08_1___RL2_n, __A08_1___WL2, __A08_1___WL2, WL02_n, GND, __A08_1___MWL2, __A08_1___RL2_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U8035(__A08_NET_298, A2XG_n, __A08_2___A1_n, __A08_NET_294, WYLOG_n, WL03_n, GND, WL02_n, WYDG_n, __A08_NET_293, __A08_2__Y1_n, CUG, __A08_2__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U8036(MONEX, __A08_NET_298, __A08_2__X1_n, CLXC, CUG, __A08_2__X1, GND, __A08_2__Y1_n, __A08_NET_294, __A08_NET_293, __A08_2__Y1, __A08_2__X1_n, __A08_2__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8037(__A08_NET_302, __A08_2__X1_n, __A08_2__Y1_n, __A08_2___XUY1, __A08_2__X1, __A08_2__Y1, GND, __A08_NET_302, __A08_2___XUY1, __A08_NET_299, __A08_NET_302, __A08_2___SUMA1, __A08_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8038( ,  , __A08_2___SUMA1, __A08_2___SUMB1, RULOG_n, __A08_NET_280, GND, __A08_NET_284, XUY05_n, __A08_2___XUY1, __A08_2___CI_IN,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U8039(__A08_2___CI_IN, __A08_NET_300, __A08_2___G1_n, __A08_2___GEM1, __A08_2___RL1_n, __A08_2___WL1, GND, WL03_n, __A08_2___WL1, __A08_2___MWL1, __A08_2___RL1_n, __A08_NET_250, __A08_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8040(__A08_2___SUMB1, __A08_NET_299, __A08_NET_300, __A08_NET_283, WAG_n, WL03_n, GND, WL05_n, WALSG_n, __A08_NET_285, __A08_2___A1_n, CAG, __A08_NET_281, VCC, SIM_RST, SIM_CLK);
    assign CO06 = CO06_U8041_2;
    assign __A08_2___RL1_n = __A08_2___RL1_n_U8041_4;
    assign __A08_2___L1_n = __A08_2___L1_n_U8041_6;
    assign __A08_2___Z1_n = __A08_2___Z1_n_U8041_8;
    assign __A08_2___RL1_n = __A08_2___RL1_n_U8041_10;
    assign __A08_2___RL1_n = __A08_2___RL1_n_U8041_12;
    U74LVC07 U8041(__A08_NET_284, CO06_U8041_2, __A08_NET_279, __A08_2___RL1_n_U8041_4, __A08_NET_291, __A08_2___L1_n_U8041_6, GND, __A08_2___Z1_n_U8041_8, __A08_NET_314, __A08_2___RL1_n_U8041_10, __A08_NET_315, __A08_2___RL1_n_U8041_12, __A08_NET_313, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U8042(__A08_NET_283, __A08_NET_285, __A08_NET_280, __A08_NET_278, CH03, __A08_NET_279, GND, __A08_NET_291, __A08_NET_282, __A08_NET_289, __A08_NET_290, __A08_2___A1_n, __A08_NET_281, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8043(__A08_NET_278, RAG_n, __A08_2___A1_n, __A08_NET_282, WLG_n, WL03_n, GND, G06_n, G2LSG_n, __A08_NET_289, __A08_2___L1_n, CLG1G, __A08_NET_290, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8044( ,  ,  ,  ,  ,  , GND, __A08_2___RL_OUT_1, RLG_n, __A08_2___L1_n, GND,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U8045( ,  ,  , __A08_NET_287, WQG_n, WL03_n, GND, __A08_NET_287, __A08_NET_286, __A08_2___Q1_n, __A08_2___Q1_n, CQG, __A08_NET_286, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U8046(__A08_NET_288, RQG_n, __A08_2___Q1_n, __A08_NET_317, WZG_n, WL03_n, GND, __A08_NET_317, __A08_NET_316, __A08_NET_314, __A08_2___Z1_n, CZG, __A08_NET_316, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U8047(__A08_NET_312, RZG_n, __A08_2___Z1_n, __A08_NET_321, WBG_n, WL03_n, GND, __A08_NET_321, __A08_NET_322, __A08_2___B1_n, __A08_2___B1_n, CBG, __A08_NET_322, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8048(__A08_NET_319, RBLG_n, __A08_2___B1_n, __A08_NET_320, __A08_NET_322, RCG_n, GND, WL02_n, WG3G_n, __A08_NET_309, WL04_n, WG4G_n, __A08_NET_308, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8049(__A08_2___RL_OUT_1, __A08_NET_288, MDT03, R1C, R15, __A08_NET_313, GND, __A08_NET_318, __A08_NET_319, __A08_NET_320, __A08_NET_305, __A08_NET_315, __A08_NET_312, VCC, SIM_RST, SIM_CLK);
    assign CO06 = CO06_U8050_2;
    assign __A08_2___RL1_n = __A08_2___RL1_n_U8050_4;
    assign __A08_2___G1_n = __A08_2___G1_n_U8050_6;
    assign __A08_2___G1_n = __A08_2___G1_n_U8050_8;
    assign __A08_2___RL2_n = __A08_2___RL2_n_U8050_10;
    assign L04_n = L04_n_U8050_12;
    U74LVC07 U8050(__A08_NET_263, CO06_U8050_2, __A08_NET_318, __A08_2___RL1_n_U8050_4, __A08_NET_304, __A08_2___G1_n_U8050_6, GND, __A08_2___G1_n_U8050_8, __A08_NET_303, __A08_2___RL2_n_U8050_10, __A08_NET_230, L04_n_U8050_12, __A08_NET_240, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8051(__A08_NET_307, L2GDG_n, L02_n, __A08_NET_306, WG1G_n, WL03_n, GND, __A08_2___G1_n, CGG, G03, RGG_n, __A08_2___G1_n, __A08_NET_305, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1, 0) U8052(__A08_NET_304, G03ED, SA03, __A08_NET_309, __A08_NET_308, __A08_NET_311, GND, __A08_NET_310, G04ED, SA04, __A08_NET_257, __A08_NET_256, __A08_NET_255, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U8053(__A08_NET_307, __A08_NET_306,  ,  ,  ,  , GND,  ,  ,  ,  , __A08_NET_303, G03, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8054(__A08_NET_251, A2XG_n, __A08_2___A2_n, __A08_NET_253, WYLOG_n, WL04_n, GND, WL03_n, WYDG_n, __A08_NET_252, __A08_2__Y2_n, CUG, __A08_2__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U8055(MONEX, __A08_NET_251, __A08_2__X2_n, CLXC, CUG, __A08_2__X2, GND, __A08_2__Y2_n, __A08_NET_253, __A08_NET_252, __A08_2__Y2, __A08_2__X2_n, __A08_2__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8056(__A08_NET_245, __A08_2__X2_n, __A08_2__Y2_n, __A08_2___XUY2, __A08_2__X2, __A08_2__Y2, GND,  ,  ,  , __A08_NET_245, __A08_2___XUY2, __A08_NET_248, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8057( ,  , __A08_NET_245, __A08_2___SUMA2, __A08_2___CO_IN, CI05_n, GND, __A08_NET_249, __A08_2___SUMA2, __A08_2___SUMB2, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U8058(__A08_2___SUMB2, __A08_NET_248, __A08_NET_250, __A08_NET_234, WAG_n, WL04_n, GND, WL06_n, WALSG_n, __A08_NET_233, __A08_2___A2_n, CAG, __A08_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U8059(__A08_NET_234, __A08_NET_233, __A08_NET_249, __A08_NET_235, CH04, __A08_NET_230, GND, __A08_NET_240, __A08_NET_268, __A08_NET_269, __A08_NET_270, __A08_2___A2_n, __A08_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8060(__A08_NET_235, RAG_n, __A08_2___A2_n, __A08_NET_268, WLG_n, WL04_n, GND, G07_n, G2LSG_n, __A08_NET_269, L04_n, CLG1G, __A08_NET_270, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8061(RLG_n, L04_n, __A08_2___RL_OUT_2, __A08_NET_236, __A08_NET_242, __A08_NET_241, GND, __A08_NET_231, MDT04, R1C, R15, __A08_2___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U8062(__A08_NET_272, WQG_n, WL04_n, __A08_2___Q2_n, __A08_NET_272, __A08_NET_271, GND, __A08_2___Q2_n, CQG, __A08_NET_271, RQG_n, __A08_2___Q2_n, __A08_NET_236, VCC, SIM_RST, SIM_CLK);
    assign __A08_2___RL2_n = __A08_2___RL2_n_U8063_2;
    assign __A08_2___Z2_n = __A08_2___Z2_n_U8063_4;
    assign __A08_2___RL2_n = __A08_2___RL2_n_U8063_6;
    assign __A08_2___RL2_n = __A08_2___RL2_n_U8063_8;
    assign __A08_2___G2_n = __A08_2___G2_n_U8063_10;
    assign __A08_2___G2_n = __A08_2___G2_n_U8063_12;
    U74LVC07 U8063(__A08_NET_241, __A08_2___RL2_n_U8063_2, __A08_NET_238, __A08_2___Z2_n_U8063_4, __A08_NET_231, __A08_2___RL2_n_U8063_6, GND, __A08_2___RL2_n_U8063_8, __A08_NET_273, __A08_2___G2_n_U8063_10, __A08_NET_255, __A08_2___G2_n_U8063_12, __A08_NET_262, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U8064(__A08_NET_237, WZG_n, WL04_n, __A08_NET_238, __A08_NET_237, __A08_NET_239, GND, __A08_2___Z2_n, CZG, __A08_NET_239, RZG_n, __A08_2___Z2_n, __A08_NET_242, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U8065(__A08_NET_276, WBG_n, WL04_n, __A08_2___B2_n, __A08_NET_276, __A08_NET_277, GND, __A08_2___B2_n, CBG, __A08_NET_277, RBLG_n, __A08_2___B2_n, __A08_NET_275, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U8066(__A08_NET_275, __A08_NET_274, __A08_NET_261, __A08_NET_260, G04, __A08_NET_262, GND,  ,  ,  ,  , __A08_NET_273, __A08_NET_254, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8067(__A08_NET_274, __A08_NET_277, RCG_n, __A08_NET_257, WL03_n, WG3G_n, GND, WL05_n, WG4G_n, __A08_NET_256, L2GDG_n, __A08_2___L1_n, __A08_NET_261, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8068(__A08_NET_260, WG1G_n, WL04_n, G04, __A08_2___G2_n, CGG, GND, RGG_n, __A08_2___G2_n, __A08_NET_254,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U8069(__A08_2___G2_n, __A08_2___GEM2, __A08_2___RL2_n, __A08_2___WL2, __A08_2___WL2, WL04_n, GND, __A08_2___MWL2, __A08_2___RL2_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC4002 U8070(__A08_1___SUMA1, __A08_NET_209, XUY01_n, CI01_n, GND, __A08_NET_174, GND, __A08_NET_173, __A08_NET_152, XUY02_n, __A08_1___CI_INTERNAL, WHOMP, __A08_1___SUMA2, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U8071(__A08_2___SUMA1, __A08_NET_302, __A08_2___XUY1, __A08_2___CI_IN, GND, __A08_NET_267, GND, __A08_NET_266, __A08_NET_245, __A08_2___XUY2, __A08_2___CI_INTERNAL, WHOMP, __A08_2___SUMA2, VCC, SIM_RST, SIM_CLK);


    U74HC02 U9001(__A09_NET_198, A2XG_n, __A09_1___A1_n, __A09_NET_193, WYLOG_n, WL05_n, GND, WL04_n, WYDG_n, __A09_NET_192, __A09_1__Y1_n, CUG, __A09_1__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U9002(MONEX, __A09_NET_198, __A09_1__X1_n, CLXC, CUG, __A09_1__X1, GND, __A09_1__Y1_n, __A09_NET_193, __A09_NET_192, __A09_1__Y1, __A09_1__X1_n, __A09_1__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9003(__A09_NET_202, __A09_1__X1_n, __A09_1__Y1_n, XUY05_n, __A09_1__X1, __A09_1__Y1, GND, __A09_NET_202, XUY05_n, __A09_NET_200, __A09_NET_202, __A09_1___SUMA1, __A09_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9004( ,  , __A09_1___SUMA1, __A09_1___SUMB1, RULOG_n, __A09_NET_180, GND, __A09_NET_184, __A09_2___XUY1, XUY05_n, CI05_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U9005(CI05_n, __A09_NET_199, G05_n, __A09_1___GEM1, __A09_1___RL1_n, __A09_1___WL1, GND, WL05_n, __A09_1___WL1, __A09_1___MWL1, __A09_1___RL1_n, __A09_NET_150, __A09_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9006(__A09_1___SUMB1, __A09_NET_200, __A09_NET_199, __A09_NET_183, WAG_n, WL05_n, GND, WL07_n, WALSG_n, __A09_NET_185, __A09_1___A1_n, CAG, __A09_NET_181, VCC, SIM_RST, SIM_CLK);
    assign __A09_2___CO_IN = __A09_2___CO_IN_U9007_2;
    assign __A09_1___RL1_n = __A09_1___RL1_n_U9007_4;
    assign __A09_1___L1_n = __A09_1___L1_n_U9007_6;
    assign __A09_1___Z1_n = __A09_1___Z1_n_U9007_8;
    assign __A09_1___RL1_n = __A09_1___RL1_n_U9007_10;
    assign __A09_1___RL1_n = __A09_1___RL1_n_U9007_12;
    U74LVC07 U9007(__A09_NET_184, __A09_2___CO_IN_U9007_2, __A09_NET_178, __A09_1___RL1_n_U9007_4, __A09_NET_191, __A09_1___L1_n_U9007_6, GND, __A09_1___Z1_n_U9007_8, __A09_NET_214, __A09_1___RL1_n_U9007_10, __A09_NET_215, __A09_1___RL1_n_U9007_12, __A09_NET_213, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9008(__A09_NET_179, RAG_n, __A09_1___A1_n, __A09_NET_182, WLG_n, WL05_n, GND, __A09_2___G2_n, G2LSG_n, __A09_NET_189, __A09_1___L1_n, CLG1G, __A09_NET_190, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U9009( ,  ,  , __A09_NET_187, WQG_n, WL05_n, GND, __A09_NET_187, __A09_NET_186, __A09_1___Q1_n, __A09_1___Q1_n, CQG, __A09_NET_186, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U9010(__A09_NET_188, RQG_n, __A09_1___Q1_n, __A09_NET_217, WZG_n, WL05_n, GND, __A09_NET_217, __A09_NET_216, __A09_NET_214, __A09_1___Z1_n, CZG, __A09_NET_216, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9011(__A09_1___RL_OUT_1, __A09_NET_188, MDT05, R1C, GND, __A09_NET_213, GND, __A09_NET_220, __A09_NET_218, __A09_NET_219, __A09_NET_205, __A09_NET_215, __A09_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U9012(__A09_NET_212, RZG_n, __A09_1___Z1_n, __A09_NET_221, WBG_n, WL05_n, GND, __A09_NET_221, __A09_NET_222, __A09_1___B1_n, __A09_1___B1_n, CBG, __A09_NET_222, VCC, SIM_RST, SIM_CLK);
    assign __A09_2___CO_IN = __A09_2___CO_IN_U9013_2;
    assign __A09_1___RL1_n = __A09_1___RL1_n_U9013_4;
    assign G05_n = G05_n_U9013_6;
    assign G05_n = G05_n_U9013_8;
    assign __A09_1___RL2_n = __A09_1___RL2_n_U9013_10;
    assign __A09_1___L2_n = __A09_1___L2_n_U9013_12;
    U74LVC07 U9013(__A09_NET_163, __A09_2___CO_IN_U9013_2, __A09_NET_220, __A09_1___RL1_n_U9013_4, __A09_NET_204, G05_n_U9013_6, GND, G05_n_U9013_8, __A09_NET_203, __A09_1___RL2_n_U9013_10, __A09_NET_130, __A09_1___L2_n_U9013_12, __A09_NET_140, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9014(__A09_NET_218, RBLG_n, __A09_1___B1_n, __A09_NET_219, __A09_NET_222, RCG_n, GND, WL04_n, WG3G_n, __A09_NET_209, WL06_n, WG4G_n, __A09_NET_208, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U9015(__A09_NET_183, __A09_NET_185, __A09_NET_180, __A09_NET_179, CH05, __A09_NET_178, GND, __A09_NET_191, __A09_NET_182, __A09_NET_189, __A09_NET_190, __A09_1___A1_n, __A09_NET_181, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9016(__A09_NET_207, L2GDG_n, L04_n, __A09_NET_206, WG1G_n, WL05_n, GND, G05_n, CGG, G05, RGG_n, G05_n, __A09_NET_205, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U9017(__A09_NET_207, __A09_NET_206, GND, __A09_2___XUY2, XUY06_n, __A09_NET_163, GND, __A09_1___RL_OUT_1, RLG_n, __A09_1___L1_n, GND, __A09_NET_203, G05, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1, 0) U9018(__A09_NET_204, G05ED, SA05, __A09_NET_209, __A09_NET_208, __A09_NET_211, GND, __A09_NET_210, G06ED, SA06, __A09_NET_157, __A09_NET_156, __A09_NET_155, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9019(__A09_NET_151, A2XG_n, __A09_1___A2_n, __A09_NET_153, WYLOG_n, WL06_n, GND, WL05_n, WYDG_n, __A09_NET_152, __A09_1__Y2_n, CUG, __A09_1__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U9020(MONEX, __A09_NET_151, __A09_1__X2_n, CLXC, CUG, __A09_1__X2, GND, __A09_1__Y2_n, __A09_NET_153, __A09_NET_152, __A09_1__Y2, __A09_1__X2_n, __A09_1__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9021(__A09_NET_145, __A09_1__X2_n, __A09_1__Y2_n, XUY06_n, __A09_1__X2, __A09_1__Y2, GND,  ,  ,  , __A09_NET_145, XUY06_n, __A09_NET_148, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9022( ,  , __A09_NET_145, __A09_1___SUMA2, CO06, __A09_2___CI_IN, GND, __A09_NET_149, __A09_1___SUMA2, __A09_1___SUMB2, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U9023(__A09_1___SUMB2, __A09_NET_148, __A09_NET_150, __A09_NET_134, WAG_n, WL06_n, GND, WL08_n, WALSG_n, __A09_NET_133, __A09_1___A2_n, CAG, __A09_NET_132, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U9024(__A09_NET_134, __A09_NET_133, __A09_NET_149, __A09_NET_135, CH06, __A09_NET_130, GND, __A09_NET_140, __A09_NET_168, __A09_NET_169, __A09_NET_170, __A09_1___A2_n, __A09_NET_132, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9025(__A09_NET_135, RAG_n, __A09_1___A2_n, __A09_NET_168, WLG_n, WL06_n, GND, G09_n, G2LSG_n, __A09_NET_169, __A09_1___L2_n, CLG1G, __A09_NET_170, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9026(RLG_n, __A09_1___L2_n, __A09_1___RL_OUT_2, __A09_NET_136, __A09_NET_142, __A09_NET_141, GND, __A09_NET_131, MDT06, R1C, GND, __A09_1___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U9027(__A09_NET_172, WQG_n, WL06_n, __A09_1___Q2_n, __A09_NET_172, __A09_NET_171, GND, __A09_1___Q2_n, CQG, __A09_NET_171, RQG_n, __A09_1___Q2_n, __A09_NET_136, VCC, SIM_RST, SIM_CLK);
    assign __A09_1___RL2_n = __A09_1___RL2_n_U9028_2;
    assign __A09_1___Z2_n = __A09_1___Z2_n_U9028_4;
    assign __A09_1___RL2_n = __A09_1___RL2_n_U9028_6;
    assign __A09_1___RL2_n = __A09_1___RL2_n_U9028_8;
    assign G06_n = G06_n_U9028_10;
    assign G06_n = G06_n_U9028_12;
    U74LVC07 U9028(__A09_NET_141, __A09_1___RL2_n_U9028_2, __A09_NET_138, __A09_1___Z2_n_U9028_4, __A09_NET_131, __A09_1___RL2_n_U9028_6, GND, __A09_1___RL2_n_U9028_8, __A09_NET_173, G06_n_U9028_10, __A09_NET_155, G06_n_U9028_12, __A09_NET_162, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U9029(__A09_NET_137, WZG_n, WL06_n, __A09_NET_138, __A09_NET_137, __A09_NET_139, GND, __A09_1___Z2_n, CZG, __A09_NET_139, RZG_n, __A09_1___Z2_n, __A09_NET_142, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U9030(__A09_NET_176, WBG_n, WL06_n, __A09_1___B2_n, __A09_NET_176, __A09_NET_177, GND, __A09_1___B2_n, CBG, __A09_NET_177, RBLG_n, __A09_1___B2_n, __A09_NET_175, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U9031(__A09_NET_175, __A09_NET_174, __A09_NET_161, __A09_NET_160, G06, __A09_NET_162, GND, __A09_NET_256, GND, XUY10_n, __A09_2___XUY2, __A09_NET_173, __A09_NET_154, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9032(__A09_NET_174, __A09_NET_177, RCG_n, __A09_NET_157, WL05_n, WG3G_n, GND, WL07_n, WG4G_n, __A09_NET_156, L2GDG_n, __A09_1___L1_n, __A09_NET_161, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9033(__A09_NET_160, WG1G_n, WL06_n, G06, G06_n, CGG, GND, RGG_n, G06_n, __A09_NET_154,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U9034(G06_n, __A09_1___GEM2, __A09_1___RL2_n, __A09_1___WL2, __A09_1___WL2, WL06_n, GND, __A09_1___MWL2, __A09_1___RL2_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U9035(__A09_NET_291, A2XG_n, __A09_2___A1_n, __A09_NET_287, WYLOG_n, WL07_n, GND, WL06_n, WYDG_n, __A09_NET_286, __A09_2__Y1_n, CUG, __A09_2__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U9036(MONEX, __A09_NET_291, __A09_2__X1_n, CLXC, CUG, __A09_2__X1, GND, __A09_2__Y1_n, __A09_NET_287, __A09_NET_286, __A09_2__Y1, __A09_2__X1_n, __A09_2__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9037(__A09_NET_295, __A09_2__X1_n, __A09_2__Y1_n, __A09_2___XUY1, __A09_2__X1, __A09_2__Y1, GND, __A09_NET_295, __A09_2___XUY1, __A09_NET_292, __A09_NET_295, __A09_2___SUMA1, __A09_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9038( ,  , __A09_2___SUMA1, __A09_2___SUMB1, RULOG_n, __A09_NET_273, GND, __A09_NET_277, XUY09_n, __A09_2___XUY1, __A09_2___CI_IN,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U9039(__A09_2___CI_IN, __A09_NET_293, G07_n, __A09_2___GEM1, __A09_2___RL1_n, __A09_2___WL1, GND, WL07_n, __A09_2___WL1, __A09_2___MWL1, __A09_2___RL1_n, __A09_NET_243, __A09_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9040(__A09_2___SUMB1, __A09_NET_292, __A09_NET_293, __A09_NET_276, WAG_n, WL07_n, GND, WL09_n, WALSG_n, __A09_NET_278, __A09_2___A1_n, CAG, __A09_NET_274, VCC, SIM_RST, SIM_CLK);
    assign CO10 = CO10_U9041_2;
    assign __A09_2___RL1_n = __A09_2___RL1_n_U9041_4;
    assign __A09_2___L1_n = __A09_2___L1_n_U9041_6;
    assign __A09_2___Z1_n = __A09_2___Z1_n_U9041_8;
    assign __A09_2___RL1_n = __A09_2___RL1_n_U9041_10;
    assign __A09_2___RL1_n = __A09_2___RL1_n_U9041_12;
    U74LVC07 U9041(__A09_NET_277, CO10_U9041_2, __A09_NET_272, __A09_2___RL1_n_U9041_4, __A09_NET_284, __A09_2___L1_n_U9041_6, GND, __A09_2___Z1_n_U9041_8, __A09_NET_307, __A09_2___RL1_n_U9041_10, __A09_NET_308, __A09_2___RL1_n_U9041_12, __A09_NET_306, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U9042(__A09_NET_276, __A09_NET_278, __A09_NET_273, __A09_NET_271, CH07, __A09_NET_272, GND, __A09_NET_284, __A09_NET_275, __A09_NET_282, __A09_NET_283, __A09_2___A1_n, __A09_NET_274, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9043(__A09_NET_271, RAG_n, __A09_2___A1_n, __A09_NET_275, WLG_n, WL07_n, GND, G10_n, G2LSG_n, __A09_NET_282, __A09_2___L1_n, CLG1G, __A09_NET_283, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9044( ,  ,  ,  ,  ,  , GND, __A09_2___RL_OUT_1, RLG_n, __A09_2___L1_n, GND,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U9045( ,  ,  , __A09_NET_280, WQG_n, WL07_n, GND, __A09_NET_280, __A09_NET_279, __A09_2___Q1_n, __A09_2___Q1_n, CQG, __A09_NET_279, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U9046(__A09_NET_281, RQG_n, __A09_2___Q1_n, __A09_NET_310, WZG_n, WL07_n, GND, __A09_NET_310, __A09_NET_309, __A09_NET_307, __A09_2___Z1_n, CZG, __A09_NET_309, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U9047(__A09_NET_305, RZG_n, __A09_2___Z1_n, __A09_NET_314, WBG_n, WL07_n, GND, __A09_NET_314, __A09_NET_315, __A09_2___B1_n, __A09_2___B1_n, CBG, __A09_NET_315, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9048(__A09_NET_312, RBLG_n, __A09_2___B1_n, __A09_NET_313, __A09_NET_315, RCG_n, GND, WL06_n, WG3G_n, __A09_NET_302, WL08_n, WG4G_n, __A09_NET_301, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9049(__A09_2___RL_OUT_1, __A09_NET_281, MDT07, R1C, GND, __A09_NET_306, GND, __A09_NET_311, __A09_NET_312, __A09_NET_313, __A09_NET_298, __A09_NET_308, __A09_NET_305, VCC, SIM_RST, SIM_CLK);
    assign CO10 = CO10_U9050_2;
    assign __A09_2___RL1_n = __A09_2___RL1_n_U9050_4;
    assign G07_n = G07_n_U9050_6;
    assign G07_n = G07_n_U9050_8;
    assign __A09_2___RL2_n = __A09_2___RL2_n_U9050_10;
    assign L08_n = L08_n_U9050_12;
    U74LVC07 U9050(__A09_NET_256, CO10_U9050_2, __A09_NET_311, __A09_2___RL1_n_U9050_4, __A09_NET_297, G07_n_U9050_6, GND, G07_n_U9050_8, __A09_NET_296, __A09_2___RL2_n_U9050_10, __A09_NET_223, L08_n_U9050_12, __A09_NET_233, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9051(__A09_NET_300, L2GDG_n, __A09_1___L2_n, __A09_NET_299, WG1G_n, WL07_n, GND, G07_n, CGG, G07, RGG_n, G07_n, __A09_NET_298, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1, 0) U9052(__A09_NET_297, G07ED, SA07, __A09_NET_302, __A09_NET_301, __A09_NET_304, GND, __A09_NET_303, GND, SA08, __A09_NET_250, __A09_NET_249, __A09_NET_248, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U9053(__A09_NET_300, __A09_NET_299,  ,  ,  ,  , GND,  ,  ,  ,  , __A09_NET_296, G07, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9054(__A09_NET_244, A2XG_n, __A09_2___A2_n, __A09_NET_246, WYLOG_n, WL08_n, GND, WL07_n, WYDG_n, __A09_NET_245, __A09_2__Y2_n, CUG, __A09_2__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U9055(MONEX, __A09_NET_244, __A09_2__X2_n, CLXC, CUG, __A09_2__X2, GND, __A09_2__Y2_n, __A09_NET_246, __A09_NET_245, __A09_2__Y2, __A09_2__X2_n, __A09_2__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9056(__A09_NET_238, __A09_2__X2_n, __A09_2__Y2_n, __A09_2___XUY2, __A09_2__X2, __A09_2__Y2, GND,  ,  ,  , __A09_NET_238, __A09_2___XUY2, __A09_NET_241, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9057( ,  , __A09_NET_238, __A09_2___SUMA2, __A09_2___CO_IN, CI09_n, GND, __A09_NET_242, __A09_2___SUMA2, __A09_2___SUMB2, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U9058(__A09_2___SUMB2, __A09_NET_241, __A09_NET_243, __A09_NET_227, WAG_n, WL08_n, GND, WL10_n, WALSG_n, __A09_NET_226, __A09_2___A2_n, CAG, __A09_NET_225, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U9059(__A09_NET_227, __A09_NET_226, __A09_NET_242, __A09_NET_228, CH08, __A09_NET_223, GND, __A09_NET_233, __A09_NET_261, __A09_NET_262, __A09_NET_263, __A09_2___A2_n, __A09_NET_225, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9060(__A09_NET_228, RAG_n, __A09_2___A2_n, __A09_NET_261, WLG_n, WL08_n, GND, G11_n, G2LSG_n, __A09_NET_262, L08_n, CLG1G, __A09_NET_263, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9061(RLG_n, L08_n, __A09_2___RL_OUT_2, __A09_NET_229, __A09_NET_235, __A09_NET_234, GND, __A09_NET_224, MDT08, R1C, GND, __A09_2___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U9062(__A09_NET_265, WQG_n, WL08_n, __A09_2___Q2_n, __A09_NET_265, __A09_NET_264, GND, __A09_2___Q2_n, CQG, __A09_NET_264, RQG_n, __A09_2___Q2_n, __A09_NET_229, VCC, SIM_RST, SIM_CLK);
    assign __A09_2___RL2_n = __A09_2___RL2_n_U9063_2;
    assign __A09_2___Z2_n = __A09_2___Z2_n_U9063_4;
    assign __A09_2___RL2_n = __A09_2___RL2_n_U9063_6;
    assign __A09_2___RL2_n = __A09_2___RL2_n_U9063_8;
    assign __A09_2___G2_n = __A09_2___G2_n_U9063_10;
    assign __A09_2___G2_n = __A09_2___G2_n_U9063_12;
    U74LVC07 U9063(__A09_NET_234, __A09_2___RL2_n_U9063_2, __A09_NET_231, __A09_2___Z2_n_U9063_4, __A09_NET_224, __A09_2___RL2_n_U9063_6, GND, __A09_2___RL2_n_U9063_8, __A09_NET_266, __A09_2___G2_n_U9063_10, __A09_NET_248, __A09_2___G2_n_U9063_12, __A09_NET_255, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U9064(__A09_NET_230, WZG_n, WL08_n, __A09_NET_231, __A09_NET_230, __A09_NET_232, GND, __A09_2___Z2_n, CZG, __A09_NET_232, RZG_n, __A09_2___Z2_n, __A09_NET_235, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U9065(__A09_NET_269, WBG_n, WL08_n, __A09_2___B2_n, __A09_NET_269, __A09_NET_270, GND, __A09_2___B2_n, CBG, __A09_NET_270, RBLG_n, __A09_2___B2_n, __A09_NET_268, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U9066(__A09_NET_268, __A09_NET_267, __A09_NET_254, __A09_NET_253, G08, __A09_NET_255, GND,  ,  ,  ,  , __A09_NET_266, __A09_NET_247, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9067(__A09_NET_267, __A09_NET_270, RCG_n, __A09_NET_250, WL07_n, WG3G_n, GND, WL09_n, WG4G_n, __A09_NET_249, L2GDG_n, __A09_2___L1_n, __A09_NET_254, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9068(__A09_NET_253, WG1G_n, WL08_n, G08, __A09_2___G2_n, CGG, GND, RGG_n, __A09_2___G2_n, __A09_NET_247,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U9069(__A09_2___G2_n, __A09_2___GEM2, __A09_2___RL2_n, __A09_2___WL2, __A09_2___WL2, WL08_n, GND, __A09_2___MWL2, __A09_2___RL2_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC4002 U9070(__A09_1___SUMA1, __A09_NET_202, XUY05_n, CI05_n, GND, __A09_NET_167, GND, __A09_NET_166, __A09_NET_145, XUY06_n, __A09_1___CI_INTERNAL, GND, __A09_1___SUMA2, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U9071(__A09_2___SUMA1, __A09_NET_295, __A09_2___XUY1, __A09_2___CI_IN, WHOMP, __A09_NET_260, GND, __A09_NET_259, __A09_NET_238, __A09_2___XUY2, __A09_2___CI_INTERNAL, GND, __A09_2___SUMA2, VCC, SIM_RST, SIM_CLK);


    U74HC02 U10001(__A10_NET_197, A2XG_n, __A10_1___A1_n, __A10_NET_192, WYLOG_n, WL09_n, GND, WL08_n, WYDG_n, __A10_NET_191, __A10_1__Y1_n, CUG, __A10_1__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U10002(MONEX, __A10_NET_197, __A10_1__X1_n, CLXC, CUG, __A10_1__X1, GND, __A10_1__Y1_n, __A10_NET_192, __A10_NET_191, __A10_1__Y1, __A10_1__X1_n, __A10_1__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10003(__A10_NET_201, __A10_1__X1_n, __A10_1__Y1_n, XUY09_n, __A10_1__X1, __A10_1__Y1, GND, __A10_NET_201, XUY09_n, __A10_NET_199, __A10_NET_201, __A10_1___SUMA1, __A10_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10004( ,  , __A10_1___SUMA1, __A10_1___SUMB1, RULOG_n, __A10_NET_179, GND, __A10_NET_183, __A10_2___XUY1, XUY09_n, CI09_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U10005(CI09_n, __A10_NET_198, G09_n, __A10_1___GEM1, __A10_1___RL1_n, __A10_1___WL1, GND, WL09_n, __A10_1___WL1, __A10_1___MWL1, __A10_1___RL1_n, __A10_NET_149, __A10_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10006(__A10_1___SUMB1, __A10_NET_199, __A10_NET_198, __A10_NET_182, WAG_n, WL09_n, GND, WL11_n, WALSG_n, __A10_NET_184, __A10_1___A1_n, CAG, __A10_NET_180, VCC, SIM_RST, SIM_CLK);
    assign __A10_2___CO_IN = __A10_2___CO_IN_U10007_2;
    assign __A10_1___RL1_n = __A10_1___RL1_n_U10007_4;
    assign __A10_1___L1_n = __A10_1___L1_n_U10007_6;
    assign __A10_1___Z1_n = __A10_1___Z1_n_U10007_8;
    assign __A10_1___RL1_n = __A10_1___RL1_n_U10007_10;
    assign __A10_1___RL1_n = __A10_1___RL1_n_U10007_12;
    U74LVC07 U10007(__A10_NET_183, __A10_2___CO_IN_U10007_2, __A10_NET_177, __A10_1___RL1_n_U10007_4, __A10_NET_190, __A10_1___L1_n_U10007_6, GND, __A10_1___Z1_n_U10007_8, __A10_NET_213, __A10_1___RL1_n_U10007_10, __A10_NET_214, __A10_1___RL1_n_U10007_12, __A10_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10008(__A10_NET_178, RAG_n, __A10_1___A1_n, __A10_NET_181, WLG_n, WL09_n, GND, __A10_2___G2_n, G2LSG_n, __A10_NET_188, __A10_1___L1_n, CLG1G, __A10_NET_189, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U10009( ,  ,  , __A10_NET_186, WQG_n, WL09_n, GND, __A10_NET_186, __A10_NET_185, __A10_1___Q1_n, __A10_1___Q1_n, CQG, __A10_NET_185, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U10010(__A10_NET_187, RQG_n, __A10_1___Q1_n, __A10_NET_216, WZG_n, WL09_n, GND, __A10_NET_216, __A10_NET_215, __A10_NET_213, __A10_1___Z1_n, CZG, __A10_NET_215, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10011(__A10_1___RL_OUT_1, __A10_NET_187, MDT09, R1C, GND, __A10_NET_212, GND, __A10_NET_219, __A10_NET_217, __A10_NET_218, __A10_NET_204, __A10_NET_214, __A10_NET_211, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U10012(__A10_NET_211, RZG_n, __A10_1___Z1_n, __A10_NET_220, WBG_n, WL09_n, GND, __A10_NET_220, __A10_NET_221, __A10_1___B1_n, __A10_1___B1_n, CBG, __A10_NET_221, VCC, SIM_RST, SIM_CLK);
    assign __A10_2___CO_IN = __A10_2___CO_IN_U10013_2;
    assign __A10_1___RL1_n = __A10_1___RL1_n_U10013_4;
    assign G09_n = G09_n_U10013_6;
    assign G09_n = G09_n_U10013_8;
    assign __A10_1___RL2_n = __A10_1___RL2_n_U10013_10;
    assign __A10_1___L2_n = __A10_1___L2_n_U10013_12;
    U74LVC07 U10013(__A10_NET_162, __A10_2___CO_IN_U10013_2, __A10_NET_219, __A10_1___RL1_n_U10013_4, __A10_NET_203, G09_n_U10013_6, GND, G09_n_U10013_8, __A10_NET_202, __A10_1___RL2_n_U10013_10, __A10_NET_129, __A10_1___L2_n_U10013_12, __A10_NET_139, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10014(__A10_NET_217, RBLG_n, __A10_1___B1_n, __A10_NET_218, __A10_NET_221, RCG_n, GND, WL08_n, WG3G_n, __A10_NET_208, WL10_n, WG4G_n, __A10_NET_207, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U10015(__A10_NET_182, __A10_NET_184, __A10_NET_179, __A10_NET_178, CH09, __A10_NET_177, GND, __A10_NET_190, __A10_NET_181, __A10_NET_188, __A10_NET_189, __A10_1___A1_n, __A10_NET_180, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10016(__A10_NET_206, L2GDG_n, L08_n, __A10_NET_205, WG1G_n, WL09_n, GND, G09_n, CGG, G09, RGG_n, G09_n, __A10_NET_204, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U10017(__A10_NET_206, __A10_NET_205, WHOMPA, __A10_2___XUY2, XUY10_n, __A10_NET_162, GND, __A10_1___RL_OUT_1, RLG_n, __A10_1___L1_n, GND, __A10_NET_202, G09, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1, 0) U10018(__A10_NET_203, GND, SA09, __A10_NET_208, __A10_NET_207, __A10_NET_210, GND, __A10_NET_209, GND, SA10, __A10_NET_156, __A10_NET_155, __A10_NET_154, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10019(__A10_NET_150, A2XG_n, __A10_1___A2_n, __A10_NET_152, WYLOG_n, WL10_n, GND, WL09_n, WYDG_n, __A10_NET_151, __A10_1__Y2_n, CUG, __A10_1__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U10020(MONEX, __A10_NET_150, __A10_1__X2_n, CLXC, CUG, __A10_1__X2, GND, __A10_1__Y2_n, __A10_NET_152, __A10_NET_151, __A10_1__Y2, __A10_1__X2_n, __A10_1__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10021(__A10_NET_144, __A10_1__X2_n, __A10_1__Y2_n, XUY10_n, __A10_1__X2, __A10_1__Y2, GND,  ,  ,  , __A10_NET_144, XUY10_n, __A10_NET_147, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10022( ,  , __A10_NET_144, __A10_1___SUMA2, CO10, __A10_2___CI_IN, GND, __A10_NET_148, __A10_1___SUMA2, __A10_1___SUMB2, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U10023(__A10_1___SUMB2, __A10_NET_147, __A10_NET_149, __A10_NET_133, WAG_n, WL10_n, GND, WL12_n, WALSG_n, __A10_NET_132, __A10_1___A2_n, CAG, __A10_NET_131, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U10024(__A10_NET_133, __A10_NET_132, __A10_NET_148, __A10_NET_134, CH10, __A10_NET_129, GND, __A10_NET_139, __A10_NET_167, __A10_NET_168, __A10_NET_169, __A10_1___A2_n, __A10_NET_131, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10025(__A10_NET_134, RAG_n, __A10_1___A2_n, __A10_NET_167, WLG_n, WL10_n, GND, G13_n, G2LSG_n, __A10_NET_168, __A10_1___L2_n, CLG1G, __A10_NET_169, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10026(RLG_n, __A10_1___L2_n, __A10_1___RL_OUT_2, __A10_NET_135, __A10_NET_141, __A10_NET_140, GND, __A10_NET_130, MDT10, R1C, GND, __A10_1___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U10027(__A10_NET_171, WQG_n, WL10_n, __A10_1___Q2_n, __A10_NET_171, __A10_NET_170, GND, __A10_1___Q2_n, CQG, __A10_NET_170, RQG_n, __A10_1___Q2_n, __A10_NET_135, VCC, SIM_RST, SIM_CLK);
    assign __A10_1___RL2_n = __A10_1___RL2_n_U10028_2;
    assign __A10_1___Z2_n = __A10_1___Z2_n_U10028_4;
    assign __A10_1___RL2_n = __A10_1___RL2_n_U10028_6;
    assign __A10_1___RL2_n = __A10_1___RL2_n_U10028_8;
    assign G10_n = G10_n_U10028_10;
    assign G10_n = G10_n_U10028_12;
    U74LVC07 U10028(__A10_NET_140, __A10_1___RL2_n_U10028_2, __A10_NET_137, __A10_1___Z2_n_U10028_4, __A10_NET_130, __A10_1___RL2_n_U10028_6, GND, __A10_1___RL2_n_U10028_8, __A10_NET_172, G10_n_U10028_10, __A10_NET_154, G10_n_U10028_12, __A10_NET_161, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U10029(__A10_NET_136, WZG_n, WL10_n, __A10_NET_137, __A10_NET_136, __A10_NET_138, GND, __A10_1___Z2_n, CZG, __A10_NET_138, RZG_n, __A10_1___Z2_n, __A10_NET_141, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U10030(__A10_NET_175, WBG_n, WL10_n, __A10_1___B2_n, __A10_NET_175, __A10_NET_176, GND, __A10_1___B2_n, CBG, __A10_NET_176, RBLG_n, __A10_1___B2_n, __A10_NET_174, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U10031(__A10_NET_174, __A10_NET_173, __A10_NET_160, __A10_NET_159, G10, __A10_NET_161, GND, __A10_NET_255, GND, XUY14_n, __A10_2___XUY2, __A10_NET_172, __A10_NET_153, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10032(__A10_NET_173, __A10_NET_176, RCG_n, __A10_NET_156, WL09_n, WG3G_n, GND, WL11_n, WG4G_n, __A10_NET_155, L2GDG_n, __A10_1___L1_n, __A10_NET_160, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10033(__A10_NET_159, WG1G_n, WL10_n, G10, G10_n, CGG, GND, RGG_n, G10_n, __A10_NET_153,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U10034(G10_n, __A10_1___GEM2, __A10_1___RL2_n, __A10_1___WL2, __A10_1___WL2, WL10_n, GND, __A10_1___MWL2, __A10_1___RL2_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U10035(__A10_NET_290, A2XG_n, __A10_2___A1_n, __A10_NET_286, WYLOG_n, WL11_n, GND, WL10_n, WYDG_n, __A10_NET_285, __A10_2__Y1_n, CUG, __A10_2__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U10036(MONEX, __A10_NET_290, __A10_2__X1_n, CLXC, CUG, __A10_2__X1, GND, __A10_2__Y1_n, __A10_NET_286, __A10_NET_285, __A10_2__Y1, __A10_2__X1_n, __A10_2__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10037(__A10_NET_294, __A10_2__X1_n, __A10_2__Y1_n, __A10_2___XUY1, __A10_2__X1, __A10_2__Y1, GND, __A10_NET_294, __A10_2___XUY1, __A10_NET_291, __A10_NET_294, __A10_2___SUMA1, __A10_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10038( ,  , __A10_2___SUMA1, __A10_2___SUMB1, RULOG_n, __A10_NET_272, GND, __A10_NET_276, XUY13_n, __A10_2___XUY1, __A10_2___CI_IN,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U10039(__A10_2___CI_IN, __A10_NET_292, G11_n, __A10_2___GEM1, __A10_2___RL1_n, __A10_2___WL1, GND, WL11_n, __A10_2___WL1, __A10_2___MWL1, __A10_2___RL1_n, __A10_NET_242, __A10_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10040(__A10_2___SUMB1, __A10_NET_291, __A10_NET_292, __A10_NET_275, WAG_n, WL11_n, GND, WL13_n, WALSG_n, __A10_NET_277, __A10_2___A1_n, CAG, __A10_NET_273, VCC, SIM_RST, SIM_CLK);
    assign CO14 = CO14_U10041_2;
    assign __A10_2___RL1_n = __A10_2___RL1_n_U10041_4;
    assign __A10_2___L1_n = __A10_2___L1_n_U10041_6;
    assign __A10_2___Z1_n = __A10_2___Z1_n_U10041_8;
    assign __A10_2___RL1_n = __A10_2___RL1_n_U10041_10;
    assign __A10_2___RL1_n = __A10_2___RL1_n_U10041_12;
    U74LVC07 U10041(__A10_NET_276, CO14_U10041_2, __A10_NET_271, __A10_2___RL1_n_U10041_4, __A10_NET_283, __A10_2___L1_n_U10041_6, GND, __A10_2___Z1_n_U10041_8, __A10_NET_306, __A10_2___RL1_n_U10041_10, __A10_NET_307, __A10_2___RL1_n_U10041_12, __A10_NET_305, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U10042(__A10_NET_275, __A10_NET_277, __A10_NET_272, __A10_NET_270, CH11, __A10_NET_271, GND, __A10_NET_283, __A10_NET_274, __A10_NET_281, __A10_NET_282, __A10_2___A1_n, __A10_NET_273, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10043(__A10_NET_270, RAG_n, __A10_2___A1_n, __A10_NET_274, WLG_n, WL11_n, GND, G14_n, G2LSG_n, __A10_NET_281, __A10_2___L1_n, CLG1G, __A10_NET_282, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10044( ,  ,  ,  ,  ,  , GND, __A10_2___RL_OUT_1, RLG_n, __A10_2___L1_n, GND,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U10045( ,  ,  , __A10_NET_279, WQG_n, WL11_n, GND, __A10_NET_279, __A10_NET_278, __A10_2___Q1_n, __A10_2___Q1_n, CQG, __A10_NET_278, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U10046(__A10_NET_280, RQG_n, __A10_2___Q1_n, __A10_NET_309, WZG_n, WL11_n, GND, __A10_NET_309, __A10_NET_308, __A10_NET_306, __A10_2___Z1_n, CZG, __A10_NET_308, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U10047(__A10_NET_304, RZG_n, __A10_2___Z1_n, __A10_NET_313, WBG_n, WL11_n, GND, __A10_NET_313, __A10_NET_314, __A10_2___B1_n, __A10_2___B1_n, CBG, __A10_NET_314, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10048(__A10_NET_311, RBHG_n, __A10_2___B1_n, __A10_NET_312, __A10_NET_314, RCG_n, GND, WL10_n, WG3G_n, __A10_NET_301, WL12_n, WG4G_n, __A10_NET_300, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10049(__A10_2___RL_OUT_1, __A10_NET_280, MDT11, R1C, GND, __A10_NET_305, GND, __A10_NET_310, __A10_NET_311, __A10_NET_312, __A10_NET_297, __A10_NET_307, __A10_NET_304, VCC, SIM_RST, SIM_CLK);
    assign CO14 = CO14_U10050_2;
    assign __A10_2___RL1_n = __A10_2___RL1_n_U10050_4;
    assign G11_n = G11_n_U10050_6;
    assign G11_n = G11_n_U10050_8;
    assign __A10_2___RL2_n = __A10_2___RL2_n_U10050_10;
    assign L12_n = L12_n_U10050_12;
    U74LVC07 U10050(__A10_NET_255, CO14_U10050_2, __A10_NET_310, __A10_2___RL1_n_U10050_4, __A10_NET_296, G11_n_U10050_6, GND, G11_n_U10050_8, __A10_NET_295, __A10_2___RL2_n_U10050_10, __A10_NET_222, L12_n_U10050_12, __A10_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10051(__A10_NET_299, L2GDG_n, __A10_1___L2_n, __A10_NET_298, WG1G_n, WL11_n, GND, G11_n, CGG, G11, RGG_n, G11_n, __A10_NET_297, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1, 0) U10052(__A10_NET_296, GND, SA11, __A10_NET_301, __A10_NET_300, __A10_NET_303, GND, __A10_NET_302, GND, SA12, __A10_NET_249, __A10_NET_248, __A10_NET_247, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U10053(__A10_NET_299, __A10_NET_298,  ,  ,  ,  , GND,  ,  ,  ,  , __A10_NET_295, G11, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10054(__A10_NET_243, A2XG_n, __A10_2___A2_n, __A10_NET_245, WYLOG_n, WL12_n, GND, WL11_n, WYDG_n, __A10_NET_244, __A10_2__Y2_n, CUG, __A10_2__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U10055(MONEX, __A10_NET_243, __A10_2__X2_n, CLXC, CUG, __A10_2__X2, GND, __A10_2__Y2_n, __A10_NET_245, __A10_NET_244, __A10_2__Y2, __A10_2__X2_n, __A10_2__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10056(__A10_NET_237, __A10_2__X2_n, __A10_2__Y2_n, __A10_2___XUY2, __A10_2__X2, __A10_2__Y2, GND,  ,  ,  , __A10_NET_237, __A10_2___XUY2, __A10_NET_240, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10057( ,  , __A10_NET_237, __A10_2___SUMA2, __A10_2___CO_IN, CI13_n, GND, __A10_NET_241, __A10_2___SUMA2, __A10_2___SUMB2, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U10058(__A10_2___SUMB2, __A10_NET_240, __A10_NET_242, __A10_NET_226, WAG_n, WL12_n, GND, WL14_n, WALSG_n, __A10_NET_225, __A10_2___A2_n, CAG, __A10_NET_224, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U10059(__A10_NET_226, __A10_NET_225, __A10_NET_241, __A10_NET_227, CH12, __A10_NET_222, GND, __A10_NET_232, __A10_NET_260, __A10_NET_261, __A10_NET_262, __A10_2___A2_n, __A10_NET_224, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10060(__A10_NET_227, RAG_n, __A10_2___A2_n, __A10_NET_260, WLG_n, WL12_n, GND, G15_n, G2LSG_n, __A10_NET_261, L12_n, CLG1G, __A10_NET_262, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10061(RLG_n, L12_n, __A10_2___RL_OUT_2, __A10_NET_228, __A10_NET_234, __A10_NET_233, GND, __A10_NET_223, MDT12, R1C, GND, __A10_2___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U10062(__A10_NET_264, WQG_n, WL12_n, __A10_2___Q2_n, __A10_NET_264, __A10_NET_263, GND, __A10_2___Q2_n, CQG, __A10_NET_263, RQG_n, __A10_2___Q2_n, __A10_NET_228, VCC, SIM_RST, SIM_CLK);
    assign __A10_2___RL2_n = __A10_2___RL2_n_U10063_2;
    assign __A10_2___Z2_n = __A10_2___Z2_n_U10063_4;
    assign __A10_2___RL2_n = __A10_2___RL2_n_U10063_6;
    assign __A10_2___RL2_n = __A10_2___RL2_n_U10063_8;
    assign __A10_2___G2_n = __A10_2___G2_n_U10063_10;
    assign __A10_2___G2_n = __A10_2___G2_n_U10063_12;
    U74LVC07 U10063(__A10_NET_233, __A10_2___RL2_n_U10063_2, __A10_NET_230, __A10_2___Z2_n_U10063_4, __A10_NET_223, __A10_2___RL2_n_U10063_6, GND, __A10_2___RL2_n_U10063_8, __A10_NET_265, __A10_2___G2_n_U10063_10, __A10_NET_247, __A10_2___G2_n_U10063_12, __A10_NET_254, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U10064(__A10_NET_229, WZG_n, WL12_n, __A10_NET_230, __A10_NET_229, __A10_NET_231, GND, __A10_2___Z2_n, CZG, __A10_NET_231, RZG_n, __A10_2___Z2_n, __A10_NET_234, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U10065(__A10_NET_268, WBG_n, WL12_n, __A10_2___B2_n, __A10_NET_268, __A10_NET_269, GND, __A10_2___B2_n, CBG, __A10_NET_269, RBHG_n, __A10_2___B2_n, __A10_NET_267, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U10066(__A10_NET_267, __A10_NET_266, __A10_NET_253, __A10_NET_252, G12, __A10_NET_254, GND,  ,  ,  ,  , __A10_NET_265, __A10_NET_246, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10067(__A10_NET_266, __A10_NET_269, RCG_n, __A10_NET_249, WL11_n, WG3G_n, GND, WL13_n, WG4G_n, __A10_NET_248, L2GDG_n, __A10_2___L1_n, __A10_NET_253, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10068(__A10_NET_252, WG1G_n, WL12_n, G12, __A10_2___G2_n, CGG, GND, RGG_n, __A10_2___G2_n, __A10_NET_246,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U10069(__A10_2___G2_n, __A10_2___GEM2, __A10_2___RL2_n, __A10_2___WL2, __A10_2___WL2, WL12_n, GND, __A10_2___MWL2, __A10_2___RL2_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC4002 U10070(__A10_1___SUMA1, __A10_NET_201, XUY09_n, CI09_n, GND, __A10_NET_166, GND, __A10_NET_165, __A10_NET_144, XUY10_n, __A10_1___CI_INTERNAL, GND, __A10_1___SUMA2, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U10071(__A10_2___SUMA1, __A10_NET_294, __A10_2___XUY1, __A10_2___CI_IN, GND, __A10_NET_259, GND, __A10_NET_258, __A10_NET_237, __A10_2___XUY2, __A10_2___CI_INTERNAL, WHOMP, __A10_2___SUMA2, VCC, SIM_RST, SIM_CLK);


    U74HC02 U11001(__A11_NET_198, A2XG_n, __A11_1___A1_n, __A11_NET_193, WYHIG_n, WL13_n, GND, WL12_n, WYDG_n, __A11_NET_192, __A11_1__Y1_n, CUG, __A11_1__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U11002(MONEX, __A11_NET_198, __A11_1__X1_n, CLXC, CUG, __A11_1__X1, GND, __A11_1__Y1_n, __A11_NET_193, __A11_NET_192, __A11_1__Y1, __A11_1__X1_n, __A11_1__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11003(__A11_NET_202, __A11_1__X1_n, __A11_1__Y1_n, XUY13_n, __A11_1__X1, __A11_1__Y1, GND, __A11_NET_202, XUY13_n, __A11_NET_200, __A11_NET_202, __A11_1___SUMA1, __A11_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11004( ,  , __A11_1___SUMA1, __A11_1___SUMB1, RULOG_n, __A11_NET_180, GND, __A11_NET_184, __A11_2___XUY1, XUY13_n, CI13_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U11005(CI13_n, __A11_NET_199, G13_n, __A11_1___GEM1, __A11_1___RL1_n, __A11_1___WL1, GND, WL13_n, __A11_1___WL1, __A11_1___MWL1, __A11_1___RL1_n, __A11_NET_150, __A11_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11006(__A11_1___SUMB1, __A11_NET_200, __A11_NET_199, __A11_NET_183, WAG_n, WL13_n, GND, WL15_n, WALSG_n, __A11_NET_185, __A11_1___A1_n, CAG, __A11_NET_181, VCC, SIM_RST, SIM_CLK);
    assign __A11_2___CO_IN = __A11_2___CO_IN_U11007_2;
    assign __A11_1___RL1_n = __A11_1___RL1_n_U11007_4;
    assign __A11_1___L1_n = __A11_1___L1_n_U11007_6;
    assign __A11_1___Z1_n = __A11_1___Z1_n_U11007_8;
    assign __A11_1___RL1_n = __A11_1___RL1_n_U11007_10;
    assign __A11_1___RL1_n = __A11_1___RL1_n_U11007_12;
    U74LVC07 U11007(__A11_NET_184, __A11_2___CO_IN_U11007_2, __A11_NET_178, __A11_1___RL1_n_U11007_4, __A11_NET_191, __A11_1___L1_n_U11007_6, GND, __A11_1___Z1_n_U11007_8, __A11_NET_214, __A11_1___RL1_n_U11007_10, __A11_NET_215, __A11_1___RL1_n_U11007_12, __A11_NET_213, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11008(__A11_NET_179, RAG_n, __A11_1___A1_n, __A11_NET_182, WLG_n, WL13_n, GND, WL01_n, WALSG_n, __A11_NET_189, __A11_1___L1_n, CLG2G, __A11_NET_190, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U11009( ,  ,  , __A11_NET_187, WQG_n, WL13_n, GND, __A11_NET_187, __A11_NET_186, __A11_1___Q1_n, __A11_1___Q1_n, CQG, __A11_NET_186, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U11010(__A11_NET_188, RQG_n, __A11_1___Q1_n, __A11_NET_217, WZG_n, WL13_n, GND, __A11_NET_217, __A11_NET_216, __A11_NET_214, __A11_1___Z1_n, CZG, __A11_NET_216, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11011(__A11_1___RL_OUT_1, __A11_NET_188, MDT13, R1C, GND, __A11_NET_213, GND, __A11_NET_220, __A11_NET_218, __A11_NET_219, __A11_NET_205, __A11_NET_215, __A11_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U11012(__A11_NET_212, RZG_n, __A11_1___Z1_n, __A11_NET_221, WBG_n, WL13_n, GND, __A11_NET_221, __A11_NET_222, __A11_1___B1_n, __A11_1___B1_n, CBG, __A11_NET_222, VCC, SIM_RST, SIM_CLK);
    assign __A11_2___CO_IN = __A11_2___CO_IN_U11013_2;
    assign __A11_1___RL1_n = __A11_1___RL1_n_U11013_4;
    assign G13_n = G13_n_U11013_6;
    assign G13_n = G13_n_U11013_8;
    assign __A11_1___RL2_n = __A11_1___RL2_n_U11013_10;
    assign __A11_1___L2_n = __A11_1___L2_n_U11013_12;
    U74LVC07 U11013(__A11_NET_163, __A11_2___CO_IN_U11013_2, __A11_NET_220, __A11_1___RL1_n_U11013_4, __A11_NET_204, G13_n_U11013_6, GND, G13_n_U11013_8, __A11_NET_203, __A11_1___RL2_n_U11013_10, __A11_NET_130, __A11_1___L2_n_U11013_12, __A11_NET_140, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11014(__A11_NET_218, RBHG_n, __A11_1___B1_n, __A11_NET_219, __A11_NET_222, RCG_n, GND, WL12_n, WG3G_n, __A11_NET_209, WL14_n, WG4G_n, __A11_NET_208, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U11015(__A11_NET_183, __A11_NET_185, __A11_NET_180, __A11_NET_179, CH13, __A11_NET_178, GND, __A11_NET_191, __A11_NET_182, __A11_NET_189, __A11_NET_190, __A11_1___A1_n, __A11_NET_181, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11016(__A11_NET_207, L2GDG_n, L12_n, __A11_NET_206, WG1G_n, WL13_n, GND, G13_n, CGG, G13, RGG_n, G13_n, __A11_NET_205, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U11017(__A11_NET_207, __A11_NET_206, GND, __A11_2___XUY2, XUY14_n, __A11_NET_163, GND, __A11_1___RL_OUT_1, RLG_n, __A11_1___L1_n, GND, __A11_NET_203, G13, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1, 0) U11018(__A11_NET_204, GND, SA13, __A11_NET_209, __A11_NET_208, __A11_NET_211, GND, __A11_NET_210, GND, SA14, __A11_NET_157, __A11_NET_156, __A11_NET_155, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11019(__A11_NET_151, A2XG_n, __A11_1___A2_n, __A11_NET_153, WYHIG_n, WL14_n, GND, WL13_n, WYDG_n, __A11_NET_152, __A11_1__Y2_n, CUG, __A11_1__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U11020(MONEX, __A11_NET_151, __A11_1__X2_n, CLXC, CUG, __A11_1__X2, GND, __A11_1__Y2_n, __A11_NET_153, __A11_NET_152, __A11_1__Y2, __A11_1__X2_n, __A11_1__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11021(__A11_NET_145, __A11_1__X2_n, __A11_1__Y2_n, XUY14_n, __A11_1__X2, __A11_1__Y2, GND,  ,  ,  , __A11_NET_145, XUY14_n, __A11_NET_148, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11022( ,  , __A11_NET_145, __A11_1___SUMA2, CO14, __A11_2___CI_IN, GND, __A11_NET_149, __A11_1___SUMA2, __A11_1___SUMB2, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U11023(__A11_1___SUMB2, __A11_NET_148, __A11_NET_150, __A11_NET_134, WAG_n, WL14_n, GND, WL16_n, WALSG_n, __A11_NET_133, __A11_1___A2_n, CAG, __A11_NET_132, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U11024(__A11_NET_134, __A11_NET_133, __A11_NET_149, __A11_NET_135, CH14, __A11_NET_130, GND, __A11_NET_140, __A11_NET_168, __A11_NET_169, __A11_NET_170, __A11_1___A2_n, __A11_NET_132, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11025(__A11_NET_135, RAG_n, __A11_1___A2_n, __A11_NET_168, WLG_n, WL14_n, GND, WL02_n, WALSG_n, __A11_NET_169, __A11_1___L2_n, CLG2G, __A11_NET_170, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11026(RLG_n, __A11_1___L2_n, __A11_1___RL_OUT_2, __A11_NET_136, __A11_NET_142, __A11_NET_141, GND, __A11_NET_131, MDT14, R1C, GND, __A11_1___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U11027(__A11_NET_172, WQG_n, WL14_n, __A11_1___Q2_n, __A11_NET_172, __A11_NET_171, GND, __A11_1___Q2_n, CQG, __A11_NET_171, RQG_n, __A11_1___Q2_n, __A11_NET_136, VCC, SIM_RST, SIM_CLK);
    assign __A11_1___RL2_n = __A11_1___RL2_n_U11028_2;
    assign __A11_1___Z2_n = __A11_1___Z2_n_U11028_4;
    assign __A11_1___RL2_n = __A11_1___RL2_n_U11028_6;
    assign __A11_1___RL2_n = __A11_1___RL2_n_U11028_8;
    assign G14_n = G14_n_U11028_10;
    assign G14_n = G14_n_U11028_12;
    U74LVC07 U11028(__A11_NET_141, __A11_1___RL2_n_U11028_2, __A11_NET_138, __A11_1___Z2_n_U11028_4, __A11_NET_131, __A11_1___RL2_n_U11028_6, GND, __A11_1___RL2_n_U11028_8, __A11_NET_173, G14_n_U11028_10, __A11_NET_155, G14_n_U11028_12, __A11_NET_162, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U11029(__A11_NET_137, WZG_n, WL14_n, __A11_NET_138, __A11_NET_137, __A11_NET_139, GND, __A11_1___Z2_n, CZG, __A11_NET_139, RZG_n, __A11_1___Z2_n, __A11_NET_142, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U11030(__A11_NET_176, WBG_n, WL14_n, __A11_1___B2_n, __A11_NET_176, __A11_NET_177, GND, __A11_1___B2_n, CBG, __A11_NET_177, RBHG_n, __A11_1___B2_n, __A11_NET_175, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U11031(__A11_NET_175, __A11_NET_174, __A11_NET_161, __A11_NET_160, G14, __A11_NET_162, GND, __A11_NET_256, GND, XUY02_n, __A11_2___XUY2, __A11_NET_173, __A11_NET_154, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11032(__A11_NET_174, __A11_NET_177, RCG_n, __A11_NET_157, WL13_n, WG3G_n, GND, WL16_n, WG4G_n, __A11_NET_156, L2GDG_n, __A11_1___L1_n, __A11_NET_161, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11033(__A11_NET_160, WG1G_n, WL14_n, G14, G14_n, CGG, GND, RGG_n, G14_n, __A11_NET_154,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U11034(G14_n, __A11_1___GEM2, __A11_1___RL2_n, __A11_1___WL2, __A11_1___WL2, WL14_n, GND, __A11_1___MWL2, __A11_1___RL2_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U11035(__A11_NET_291, A2XG_n, __A11_2___A1_n, __A11_NET_287, WYHIG_n, WL15_n, GND, WL14_n, WYDG_n, __A11_NET_286, __A11_2__Y1_n, CUG, __A11_2__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U11036(BXVX, __A11_NET_291, __A11_2__X1_n, CLXC, CUG, __A11_2__X1, GND, __A11_2__Y1_n, __A11_NET_287, __A11_NET_286, __A11_2__Y1, __A11_2__X1_n, __A11_2__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11037(__A11_NET_295, __A11_2__X1_n, __A11_2__Y1_n, __A11_2___XUY1, __A11_2__X1, __A11_2__Y1, GND, __A11_NET_295, __A11_2___XUY1, __A11_NET_292, __A11_NET_295, SUMA15_n, __A11_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11038( ,  , SUMA15_n, SUMB15_n, RULOG_n, __A11_NET_273, GND, __A11_NET_277, XUY01_n, __A11_2___XUY1, __A11_2___CI_IN,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U11039(__A11_2___CI_IN, __A11_NET_293, G15_n, __A11_2___GEM1, __A11_2___RL1_n, WL15, GND, WL15_n, WL15, __A11_2___MWL1, __A11_2___RL1_n, __A11_NET_243, __A11_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11040(SUMB15_n, __A11_NET_292, __A11_NET_293, __A11_NET_276, WAG_n, WL15_n, GND, G16SW_n, WALSG_n, __A11_NET_278, __A11_2___A1_n, CAG, __A11_NET_274, VCC, SIM_RST, SIM_CLK);
    assign __A11_2___CO_OUT = __A11_2___CO_OUT_U11041_2;
    assign __A11_2___RL1_n = __A11_2___RL1_n_U11041_4;
    assign L15_n = L15_n_U11041_6;
    assign __A11_2___Z1_n = __A11_2___Z1_n_U11041_8;
    assign __A11_2___RL1_n = __A11_2___RL1_n_U11041_10;
    assign __A11_2___RL1_n = __A11_2___RL1_n_U11041_12;
    U74LVC07 U11041(__A11_NET_277, __A11_2___CO_OUT_U11041_2, __A11_NET_272, __A11_2___RL1_n_U11041_4, __A11_NET_284, L15_n_U11041_6, GND, __A11_2___Z1_n_U11041_8, __A11_NET_307, __A11_2___RL1_n_U11041_10, __A11_NET_308, __A11_2___RL1_n_U11041_12, __A11_NET_306, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U11042(__A11_NET_276, __A11_NET_278, __A11_NET_273, __A11_NET_271, CH16, __A11_NET_272, GND, __A11_NET_284, __A11_NET_275, __A11_NET_282, __A11_NET_283, __A11_2___A1_n, __A11_NET_274, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11043(__A11_NET_271, RAG_n, __A11_2___A1_n, __A11_NET_275, WLG_n, WL15_n, GND, G01_n, G2LSG_n, __A11_NET_282, L15_n, CLG1G, __A11_NET_283, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11044( ,  ,  ,  ,  ,  , GND, __A11_2___RL_OUT_1, RLG_n, L15_n, VCC,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U11045( ,  ,  , __A11_NET_280, WQG_n, WL15_n, GND, __A11_NET_280, __A11_NET_279, __A11_2___Q1_n, __A11_2___Q1_n, CQG, __A11_NET_279, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U11046(__A11_NET_281, RQG_n, __A11_2___Q1_n, __A11_NET_310, WZG_n, WL15_n, GND, __A11_NET_310, __A11_NET_309, __A11_NET_307, __A11_2___Z1_n, CZG, __A11_NET_309, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U11047(__A11_NET_305, RZG_n, __A11_2___Z1_n, __A11_NET_314, WBG_n, WL15_n, GND, __A11_NET_314, __A11_NET_315, __A11_2___B1_n, __A11_2___B1_n, CBG, __A11_NET_315, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11048(__A11_NET_312, RBHG_n, __A11_2___B1_n, __A11_NET_313, __A11_NET_315, RCG_n, GND, GND, VCC, __A11_NET_302, GND, VCC, __A11_NET_301, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11049(__A11_2___RL_OUT_1, __A11_NET_281, MDT15, R1C, __A11_2___RL_OUT_2, __A11_NET_306, GND, __A11_NET_311, __A11_NET_312, __A11_NET_313, __A11_NET_298, __A11_NET_308, __A11_NET_305, VCC, SIM_RST, SIM_CLK);
    assign __A11_2___CO_OUT = __A11_2___CO_OUT_U11050_2;
    assign __A11_2___RL1_n = __A11_2___RL1_n_U11050_4;
    assign G15_n = G15_n_U11050_6;
    assign G15_n = G15_n_U11050_8;
    assign __A11_2___RL2_n = __A11_2___RL2_n_U11050_10;
    assign __A11_2___L2_n = __A11_2___L2_n_U11050_12;
    U74LVC07 U11050(__A11_NET_256, __A11_2___CO_OUT_U11050_2, __A11_NET_311, __A11_2___RL1_n_U11050_4, __A11_NET_297, G15_n_U11050_6, GND, G15_n_U11050_8, __A11_NET_296, __A11_2___RL2_n_U11050_10, __A11_NET_223, __A11_2___L2_n_U11050_12, __A11_NET_233, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11051(__A11_NET_300, L2GDG_n, __A11_1___L2_n, __A11_NET_299, WG1G_n, WL15_n, GND, G15_n, CGG, G15, RGG_n, G15_n, __A11_NET_298, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1, 0) U11052(__A11_NET_297, GND, SA16, __A11_NET_302, __A11_NET_301, __A11_NET_304, GND, __A11_NET_303, GND, SA16, __A11_NET_250, __A11_NET_249, __A11_NET_248, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U11053(__A11_NET_300, __A11_NET_299,  ,  ,  ,  , GND,  ,  ,  ,  , __A11_NET_296, G15, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11054(__A11_NET_244, A2XG_n, __A11_2___A2_n, __A11_NET_246, WYHIG_n, WL16_n, GND, WL16_n, WYDG_n, __A11_NET_245, __A11_2__Y2_n, CUG, __A11_2__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U11055(MONEX, __A11_NET_244, __A11_2__X2_n, CLXC, CUG, __A11_2__X2, GND, __A11_2__Y2_n, __A11_NET_246, __A11_NET_245, __A11_2__Y2, __A11_2__X2_n, __A11_2__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11056(__A11_NET_238, __A11_2__X2_n, __A11_2__Y2_n, __A11_2___XUY2, __A11_2__X2, __A11_2__Y2, GND,  ,  ,  , __A11_NET_238, __A11_2___XUY2, __A11_NET_241, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11057( ,  , __A11_NET_238, SUMA16_n, __A11_2___CO_IN, EAC_n, GND, __A11_NET_242, SUMA16_n, SUMB16_n, RUG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U11058(SUMB16_n, __A11_NET_241, __A11_NET_243, __A11_NET_227, WAG_n, WL16_n, GND, G16SW_n, WALSG_n, __A11_NET_226, __A11_2___A2_n, CAG, __A11_NET_225, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 1) U11059(__A11_NET_227, __A11_NET_226, __A11_NET_242, __A11_NET_228, CH16, __A11_NET_223, GND, __A11_NET_233, __A11_NET_261, __A11_NET_262, __A11_NET_263, __A11_2___A2_n, __A11_NET_225, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11060(__A11_NET_228, RAG_n, __A11_2___A2_n, __A11_NET_261, WLG_n, WL16_n, GND, __A11_2___G2_n, G2LSG_n, __A11_NET_262, __A11_2___L2_n, CLG1G, __A11_NET_263, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11061(RLG_n, __A11_2___L2_n, __A11_2___RL_OUT_2, __A11_NET_229, __A11_NET_235, __A11_NET_234, GND, __A11_NET_224, MDT16, R1C, US2SG, __A11_2___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U11062(__A11_NET_265, WQG_n, WL16_n, __A11_2___Q2_n, __A11_NET_265, __A11_NET_264, GND, __A11_2___Q2_n, CQG, __A11_NET_264, RQG_n, __A11_2___Q2_n, __A11_NET_229, VCC, SIM_RST, SIM_CLK);
    assign __A11_2___RL2_n = __A11_2___RL2_n_U11063_2;
    assign __A11_2___Z2_n = __A11_2___Z2_n_U11063_4;
    assign __A11_2___RL2_n = __A11_2___RL2_n_U11063_6;
    assign __A11_2___RL2_n = __A11_2___RL2_n_U11063_8;
    assign __A11_2___G2_n = __A11_2___G2_n_U11063_10;
    assign __A11_2___G2_n = __A11_2___G2_n_U11063_12;
    U74LVC07 U11063(__A11_NET_234, __A11_2___RL2_n_U11063_2, __A11_NET_231, __A11_2___Z2_n_U11063_4, __A11_NET_224, __A11_2___RL2_n_U11063_6, GND, __A11_2___RL2_n_U11063_8, __A11_NET_266, __A11_2___G2_n_U11063_10, __A11_NET_248, __A11_2___G2_n_U11063_12, __A11_NET_255, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U11064(__A11_NET_230, WZG_n, WL16_n, __A11_NET_231, __A11_NET_230, __A11_NET_232, GND, __A11_2___Z2_n, CZG, __A11_NET_232, RZG_n, __A11_2___Z2_n, __A11_NET_235, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U11065(__A11_NET_269, WBG_n, WL16_n, __A11_2___B2_n, __A11_NET_269, __A11_NET_270, GND, __A11_2___B2_n, CBG, __A11_NET_270, RBHG_n, __A11_2___B2_n, __A11_NET_268, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U11066(__A11_NET_268, __A11_NET_267, __A11_NET_254, __A11_NET_253, G16, __A11_NET_255, GND,  ,  ,  ,  , __A11_NET_266, __A11_NET_247, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11067(__A11_NET_267, __A11_NET_270, RCG_n, __A11_NET_250, WL14_n, WG3G_n, GND, WL01_n, WG5G_n, __A11_NET_249, L2GDG_n, __A11_2___L2_n, __A11_NET_254, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11068(__A11_NET_253, WG2G_n, WL16_n, G16, __A11_2___G2_n, CGG, GND, RGG_n, __A11_2___G2_n, __A11_NET_247,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U11069(__A11_2___G2_n, __A11_2___GEM2, __A11_2___RL2_n, WL16, WL16, WL16_n, GND, __A11_2___MWL2, __A11_2___RL2_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC4002 U11070(__A11_1___SUMA1, __A11_NET_202, XUY13_n, CI13_n, GND, __A11_NET_167, GND, __A11_NET_166, __A11_NET_145, XUY14_n, __A11_1___CI_INTERNAL, GND, __A11_1___SUMA2, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U11071(SUMA15_n, __A11_NET_295, __A11_2___XUY1, __A11_2___CI_IN, GND, __A11_NET_260, GND, __A11_NET_259, __A11_NET_238, __A11_2___XUY2, __A11_2___CI_INTERNAL, WHOMPA, SUMA16_n, VCC, SIM_RST, SIM_CLK);


    U74HC04 U12001(G01, __A12_1__G01A_n, G02, __A12_1__G02_n, G03, __A12_1__G03_n, GND, __A12_1__PA03_n, __A12_1__PA03, __A12_NET_196, G04, __A12_NET_190, G05, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12002(G01, G02, G01, __A12_1__G02_n, __A12_1__G03_n, __A12_NET_182, GND, __A12_NET_181, __A12_1__G01A_n, G02, __A12_1__G03_n, __A12_NET_177, G03, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12003(__A12_1__G01A_n, __A12_1__G02_n, G04, G05, G06, __A12_NET_183, GND, __A12_NET_186, G04, __A12_NET_190, __A12_NET_195, __A12_NET_180, G03, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U12004(__A12_1__PA03, __A12_NET_177, __A12_NET_182, __A12_NET_181, __A12_NET_180, __A12_NET_179, GND, __A12_NET_178, __A12_NET_183, __A12_NET_186, __A12_NET_185, __A12_NET_184, __A12_1__PA06, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12005(G06, __A12_NET_195, __A12_NET_183, __A12_NET_133, __A12_1__PA06, __A12_1__PA06_n, GND, __A12_NET_189, G07, __A12_NET_127, G08, __A12_NET_174, G09, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12006(__A12_NET_196, G05, __A12_NET_196, __A12_NET_190, G06, __A12_NET_184, GND, __A12_NET_123, G07, G08, G09, __A12_NET_185, __A12_NET_195, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12007(G07, __A12_NET_127, __A12_NET_189, G08, __A12_NET_174, __A12_NET_126, GND, __A12_NET_125, __A12_NET_189, __A12_NET_127, G09, __A12_NET_122, __A12_NET_174, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U12008(__A12_1__PA09, __A12_NET_123, __A12_NET_122, __A12_NET_126, __A12_NET_125, __A12_NET_173, GND, __A12_NET_172, __A12_NET_136, __A12_NET_135, __A12_NET_138, __A12_NET_137, __A12_1__PA12, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12009(__A12_NET_123, __A12_NET_132, __A12_1__PA09, __A12_1__PA09_n, G10, __A12_NET_120, GND, __A12_NET_124, G11, __A12_NET_121, G12, __A12_NET_114, __A12_NET_136, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12010(G10, G11, G10, __A12_NET_124, __A12_NET_121, __A12_NET_135, GND, __A12_NET_138, __A12_NET_120, G11, __A12_NET_121, __A12_NET_136, G12, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12011(__A12_NET_120, __A12_NET_124, G13, G14, G16, __A12_NET_134, GND, __A12_NET_130, G13, __A12_NET_131, __A12_NET_139, __A12_NET_137, G12, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12012(__A12_1__PA12, __A12_1__PA12_n, G13, __A12_NET_140, G14, __A12_NET_131, GND, __A12_NET_139, G16, __A12_NET_113, __A12_NET_134, __A12_1__PA15_n, __A12_1__PA15, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12013(__A12_NET_140, G14, __A12_NET_140, __A12_NET_131, G16, __A12_NET_128, GND, __A12_NET_198, __A12_NET_133, __A12_NET_132, __A12_NET_114, __A12_NET_129, __A12_NET_139, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(0, 1) U12014(__A12_1__PA15, __A12_NET_134, __A12_NET_130, __A12_NET_129, __A12_NET_128, __A12_NET_200, GND, __A12_NET_199, EXTPLS, RELPLS, INHPLS, __A12_NET_118, __A12_NET_119, VCC, SIM_RST, SIM_CLK);
    U74HC02 U12015(__A12_NET_197, __A12_NET_113, G15, __A12_NET_110, TSUDO_n, __A12_1__T7PHS4_n, GND, __A12_1__G02_n, G03, __A12_NET_192, G02, __A12_1__G03_n, __A12_NET_191, VCC, SIM_RST, SIM_CLK);
    assign __A12_1__GNZRO = __A12_1__GNZRO_U12016_2;
    assign __A12_1__GNZRO = __A12_1__GNZRO_U12016_4;
    assign RELPLS = RELPLS_U12016_6;
    assign RELPLS = RELPLS_U12016_8;
    assign INHPLS = INHPLS_U12016_10;
    assign INHPLS = INHPLS_U12016_12;
    U74LVC07 U12016(__A12_NET_198, __A12_1__GNZRO_U12016_2, __A12_NET_197, __A12_1__GNZRO_U12016_4, __A12_NET_193, RELPLS_U12016_6, GND, RELPLS_U12016_8, __A12_NET_192, INHPLS_U12016_10, __A12_NET_194, INHPLS_U12016_12, __A12_NET_191, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12017(__A12_1__GNZRO, __A12_NET_109, __A12_NET_182, __A12_NET_112, __A12_NET_110, __A12_NET_111, GND, GEQZRO_n, __A12_NET_108, __A12_NET_116, RAD, __A12_1__PB09_n, __A12_1__PB09, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12018(__A12_NET_112, __A12_NET_109, __A12_NET_109, __A12_NET_111, __A12_1__G01A_n, __A12_NET_193, GND, __A12_NET_194, __A12_NET_109, G01, __A12_NET_111, EXTPLS, __A12_NET_111, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U12019(__A12_NET_108, __A12_NET_109, G02, G01, G03, __A12_NET_107, GND, __A12_NET_106, __A12_NET_151, __A12_NET_150, __A12_NET_149, __A12_NET_165, __A12_1__PB09, VCC, SIM_RST, SIM_CLK);
    U74HC02 U12020(__A12_NET_118, __A12_NET_119, T12A, RADRZ, __A12_NET_119, __A12_NET_116, GND, __A12_NET_116, __A12_NET_118, RADRG, __A12_1__PA12, __A12_1__PA15, __A12_NET_156, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12021(__A12_1__PA03, __A12_1__PA06, __A12_1__PA03, __A12_1__PA06_n, __A12_1__PA09_n, __A12_NET_150, GND, __A12_NET_149, __A12_1__PA03_n, __A12_1__PA06, __A12_1__PA09_n, __A12_NET_151, __A12_1__PA09, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(0, 1, 0) U12022(__A12_1__PA03_n, __A12_1__PA06_n, __A12_NET_142, MONPAR, SAP, __A12_NET_143, GND, __A12_NET_148, SCAD, __A12_NET_141, GOJAM, __A12_NET_165, __A12_1__PA09, VCC, SIM_RST, SIM_CLK);
    U74HC02 U12023(__A12_NET_155, __A12_1__PA12_n, __A12_1__PA15_n, __A12_1__PB15, __A12_NET_156, __A12_NET_155, GND, __A12_1__PB09_n, __A12_1__PB15, __A12_NET_166, __A12_1__PB09, __A12_1__PB15_n, __A12_NET_168, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12024(__A12_1__PB15, __A12_1__PB15_n, __A12_1__PC15, __A12_1__PC15_n, __A12_1__PC15, __A12_1__MGP_n, GND, __A12_1__GEMP, __A12_1__PC15_n, __A12_1__MSP, __A12_NET_143, __A12_1__MPAL, __A12_1__PALE, VCC, SIM_RST, SIM_CLK);
    U74HC02 U12025(__A12_1__PC15, __A12_NET_166, __A12_NET_168, __A12_NET_142, CGG, __A12_NET_143, GND, __A12_1__PC15, __A12_NET_142, __A12_NET_141, __A12_1__PC15_n, __A12_NET_143, __A12_NET_146, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12026(TPARG_n, n8XP5, T07_n, PHS4_n, FUTEXT, __A12_1__T7PHS4, GND, __A12_NET_243, XB0_n, T02_n, __A12_NET_242, __A12_NET_147, __A12_NET_146, VCC, SIM_RST, SIM_CLK);
    assign __A12_1__PALE = __A12_1__PALE_U12027_2;
    assign __A12_1__PALE = __A12_1__PALE_U12027_4;
    U74LVC07 U12027(__A12_NET_148, __A12_1__PALE_U12027_2, __A12_NET_147, __A12_1__PALE_U12027_4,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U12028(G01ED, WEDOPG_n, WL08_n, __A12_NET_233, WL08_n, WSG_n, GND, __A12_NET_233, __A12_NET_232, __A12_NET_231, __A12_NET_231, CSG, __A12_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12029(__A12_NET_231, __A12_2__S08, __A12_NET_232, __A12_2__S08_n, __A12_NET_226, __A12_2__S09, GND, __A12_2__S09_n, __A12_NET_225, __A12_2__S10, __A12_NET_229, __A12_2__S10_n, __A12_NET_228, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U12030(G02ED, WEDOPG_n, WL09_n, __A12_NET_227, WL09_n, WSG_n, GND, __A12_NET_227, __A12_NET_225, __A12_NET_226, __A12_NET_226, CSG, __A12_NET_225, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U12031(G03ED, WEDOPG_n, WL10_n, __A12_NET_230, WL10_n, WSG_n, GND, __A12_NET_230, __A12_NET_228, __A12_NET_229, __A12_NET_229, CSG, __A12_NET_228, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U12032(G04ED, WEDOPG_n, WL11_n, __A12_NET_239, WL11_n, WSG_n, GND, __A12_NET_239, __A12_NET_237, __A12_NET_238, __A12_NET_238, CSG, __A12_NET_237, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12033(__A12_NET_238, S11, __A12_NET_237, __A12_2__S11_n, __A12_NET_235, S12, GND, __A12_2__S12_n, __A12_NET_236, __A12_2__S01, __A12_NET_213, __A12_2__S01_n, __A12_NET_211, VCC, SIM_RST, SIM_CLK);
    U74HC02 U12034(G05ED, WEDOPG_n, WL12_n, __A12_NET_234, WL12_n, WSG_n, GND, EDOP_n, T12A, __A12_NET_250, __A12_NET_235, CSG, __A12_NET_236, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 0, 1) U12035(G06ED, WEDOPG_n, WL13_n, G07ED, WEDOPG_n, WL14_n, GND, WL01_n, WSG_n, __A12_NET_212, __A12_NET_212, __A12_NET_211, __A12_NET_213, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U12036(__A12_NET_211, __A12_NET_213, CSG, __A12_NET_206, WL02_n, WSG_n, GND, __A12_NET_206, __A12_NET_205, __A12_NET_204, __A12_NET_204, CSG, __A12_NET_205, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12037(__A12_NET_204, __A12_2__S02, __A12_NET_205, __A12_2__S02_n, __A12_NET_209, __A12_2__S03, GND, __A12_2__S03_n, __A12_NET_208, __A12_2__S04, __A12_NET_220, __A12_2__S04_n, __A12_NET_222, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U12038(__A12_NET_207, WL03_n, WSG_n, __A12_NET_209, __A12_NET_207, __A12_NET_208, GND, __A12_NET_209, CSG, __A12_NET_208, WL04_n, WSG_n, __A12_NET_210, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1, 0, 0, 1) U12039(__A12_NET_220, __A12_NET_210, __A12_NET_222, __A12_NET_222, __A12_NET_220, CSG, GND, WL05_n, WSG_n, __A12_NET_223, __A12_NET_223, __A12_NET_219, __A12_NET_221, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 0, 1, 0) U12040(__A12_NET_219, __A12_NET_221, CSG, __A12_NET_224, WL06_n, WSG_n, GND, __A12_NET_224, __A12_NET_217, __A12_NET_218, __A12_NET_218, __A12_NET_252, __A12_NET_217, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12041(__A12_NET_221, __A12_2__S05, __A12_NET_219, __A12_2__S05_n, __A12_NET_218, __A12_2__S06, GND, __A12_2__S06_n, __A12_NET_217, __A12_2__S07, __A12_NET_216, __A12_2__S07_n, __A12_NET_214, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 0) U12042(__A12_NET_215, WL07_n, WSG_n, __A12_NET_216, __A12_NET_215, __A12_NET_214, GND, __A12_NET_216, CSG, __A12_NET_214,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U12043(__A12_1__T7PHS4, __A12_1__T7PHS4_n,  ,  , OCTAD2, __A12_NET_242, GND, GINH, __A12_NET_249,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC4002 U12044( ,  ,  ,  ,  , __A12_NET_247, GND, __A12_NET_248, __A12_NET_244, __A12_NET_246, __A12_NET_245, __A12_NET_250, __A12_NET_249, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 1) U12046( ,  ,  , CYR_n, __A12_NET_243, __A12_NET_244, GND, CYR_n, T12A, __A12_NET_244, __A12_NET_240, __A12_NET_246, SR_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12047(__A12_NET_242, T02_n, __A12_NET_242, T02_n, XB2_n, __A12_NET_241, GND, __A12_NET_251, __A12_NET_242, T02_n, XB3_n, __A12_NET_240, XB1_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(0, 1, 0, 1) U12048(__A12_NET_246, SR_n, T12A, CYL_n, __A12_NET_241, __A12_NET_245, GND, CYL_n, T12A, __A12_NET_245, __A12_NET_251, __A12_NET_250, EDOP_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1, 0, 0) U12049(n8XP5, __A12_NET_234,  ,  ,  ,  , GND,  ,  ,  ,  , __A12_NET_235, __A12_NET_236, VCC, SIM_RST, SIM_CLK);
endmodule
