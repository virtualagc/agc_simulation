`timescale 1ns/1ps
`default_nettype none

module inout_i(VCC, GND, SIM_RST, SIM_CLK, GOJAM, CCHG_n, WCHG_n, CCH11, RCH11_n, WCH11_n, FLASH, FLASH_n, XT0_n, XT1_n, XB2_n, XB5_n, XB6_n, CHWL01_n, CHWL02_n, CHWL03_n, CHWL04_n, CHWL05_n, CHWL06_n, CHWL07_n, CHWL08_n, CHWL09_n, CHWL10_n, CHWL11_n, CHWL12_n, CHWL13_n, CHWL14_n, CH0705, CH0706, CH0707, CH1501, CH1502, CH1503, CH1504, CH3201, CH3202, CH3203, CH3204, CH3205, CH3206, CH3207, CH3208, CCH12, RCH12_n, WCH12_n, TMPOUT, CH1213, CH1214, CH1208, CH1209, CH1210, CH1211, CH1212, CHOR01_n, CHOR02_n, CHOR03_n, CHOR04_n, CHOR05_n, CHOR06_n, CHOR07_n, CHOR08_n);
    input wire VCC;
    input wire GND;
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire CCH11;
    output wire CCH12;
    input wire CCHG_n;
    input wire CH0705;
    input wire CH0706;
    input wire CH0707;
    output wire CH1208;
    output wire CH1209;
    output wire CH1210;
    output wire CH1211;
    output wire CH1212;
    output wire CH1213;
    output wire CH1214;
    input wire CH1501;
    input wire CH1502;
    input wire CH1503;
    input wire CH1504;
    input wire CH3201;
    input wire CH3202;
    input wire CH3203;
    input wire CH3204;
    input wire CH3205;
    input wire CH3206;
    input wire CH3207;
    input wire CH3208;
    output wire CHOR01_n; //FPGA#wand
    output wire CHOR02_n; //FPGA#wand
    output wire CHOR03_n; //FPGA#wand
    output wire CHOR04_n; //FPGA#wand
    output wire CHOR05_n; //FPGA#wand
    output wire CHOR06_n; //FPGA#wand
    output wire CHOR07_n; //FPGA#wand
    output wire CHOR08_n; //FPGA#wand
    input wire CHWL01_n;
    input wire CHWL02_n;
    input wire CHWL03_n;
    input wire CHWL04_n;
    input wire CHWL05_n;
    input wire CHWL06_n;
    input wire CHWL07_n;
    input wire CHWL08_n;
    input wire CHWL09_n;
    input wire CHWL10_n;
    input wire CHWL11_n;
    input wire CHWL12_n;
    input wire CHWL13_n;
    input wire CHWL14_n;
    input wire FLASH;
    input wire FLASH_n;
    input wire GOJAM;
    input wire RCH11_n;
    output wire RCH12_n;
    output wire TMPOUT;
    input wire WCH11_n;
    output wire WCH12_n;
    input wire WCHG_n;
    input wire XB2_n;
    input wire XB5_n;
    input wire XB6_n;
    input wire XT0_n;
    input wire XT1_n;
    wire __A16_1__CCH05;
    wire __A16_1__CCH06;
    wire __A16_1__CH1207;
    wire __A16_1__OT1207;
    wire __A16_1__OT1207_n;
    wire __A16_1__RCH05_n;
    wire __A16_1__RCH06_n;
    wire __A16_1__RCmXmP;
    wire __A16_1__RCmXmY;
    wire __A16_1__RCmXpP;
    wire __A16_1__RCmXpY;
    wire __A16_1__RCmYmR;
    wire __A16_1__RCmYpR;
    wire __A16_1__RCmZmR;
    wire __A16_1__RCmZpR;
    wire __A16_1__RCpXmP;
    wire __A16_1__RCpXmY;
    wire __A16_1__RCpXpP;
    wire __A16_1__RCpXpY;
    wire __A16_1__RCpYmR;
    wire __A16_1__RCpYpR;
    wire __A16_1__RCpZmR;
    wire __A16_1__RCpZpR;
    wire __A16_1__TVCNAB;
    wire __A16_1__WCH05_n;
    wire __A16_1__WCH06_n;
    wire __A16_2__COARSE;
    wire __A16_2__COMACT;
    wire __A16_2__DISDAC;
    wire __A16_2__ENERIM;
    wire __A16_2__ENEROP;
    wire __A16_2__KYRLS;
    wire __A16_2__MROLGT;
    wire __A16_2__OPEROR;
    wire __A16_2__S4BOFF;
    wire __A16_2__S4BSEQ;
    wire __A16_2__S4BTAK;
    wire __A16_2__STARON;
    wire __A16_2__UPLACT;
    wire __A16_2__VNFLSH;
    wire __A16_2__ZEROPT;
    wire __A16_2__ZIMCDU;
    wire __A16_2__ZOPCDU;
    wire __A16_NET_101;
    wire __A16_NET_102;
    wire __A16_NET_103;
    wire __A16_NET_104;
    wire __A16_NET_105;
    wire __A16_NET_106;
    wire __A16_NET_107;
    wire __A16_NET_108;
    wire __A16_NET_109;
    wire __A16_NET_110;
    wire __A16_NET_111;
    wire __A16_NET_112;
    wire __A16_NET_113;
    wire __A16_NET_114;
    wire __A16_NET_115;
    wire __A16_NET_116;
    wire __A16_NET_117;
    wire __A16_NET_118;
    wire __A16_NET_119;
    wire __A16_NET_120;
    wire __A16_NET_121;
    wire __A16_NET_122;
    wire __A16_NET_123;
    wire __A16_NET_124;
    wire __A16_NET_125;
    wire __A16_NET_126;
    wire __A16_NET_127;
    wire __A16_NET_128;
    wire __A16_NET_129;
    wire __A16_NET_130;
    wire __A16_NET_131;
    wire __A16_NET_132;
    wire __A16_NET_133;
    wire __A16_NET_134;
    wire __A16_NET_135;
    wire __A16_NET_136;
    wire __A16_NET_137;
    wire __A16_NET_138;
    wire __A16_NET_139;
    wire __A16_NET_140;
    wire __A16_NET_141;
    wire __A16_NET_142;
    wire __A16_NET_143;
    wire __A16_NET_144;
    wire __A16_NET_145;
    wire __A16_NET_146;
    wire __A16_NET_147;
    wire __A16_NET_148;
    wire __A16_NET_149;
    wire __A16_NET_150;
    wire __A16_NET_151;
    wire __A16_NET_152;
    wire __A16_NET_153;
    wire __A16_NET_154;
    wire __A16_NET_155;
    wire __A16_NET_156;
    wire __A16_NET_161;
    wire __A16_NET_162;
    wire __A16_NET_163;
    wire __A16_NET_164;
    wire __A16_NET_165;
    wire __A16_NET_168;
    wire __A16_NET_169;
    wire __A16_NET_170;
    wire __A16_NET_171;
    wire __A16_NET_172;
    wire __A16_NET_173;
    wire __A16_NET_174;
    wire __A16_NET_175;
    wire __A16_NET_176;
    wire __A16_NET_177;
    wire __A16_NET_178;
    wire __A16_NET_179;
    wire __A16_NET_180;
    wire __A16_NET_181;
    wire __A16_NET_182;
    wire __A16_NET_183;
    wire __A16_NET_184;
    wire __A16_NET_185;
    wire __A16_NET_186;
    wire __A16_NET_187;
    wire __A16_NET_188;
    wire __A16_NET_189;
    wire __A16_NET_190;
    wire __A16_NET_191;
    wire __A16_NET_192;
    wire __A16_NET_193;
    wire __A16_NET_194;
    wire __A16_NET_195;
    wire __A16_NET_196;
    wire __A16_NET_197;
    wire __A16_NET_198;
    wire __A16_NET_199;
    wire __A16_NET_200;
    wire __A16_NET_201;
    wire __A16_NET_202;
    wire __A16_NET_203;
    wire __A16_NET_204;
    wire __A16_NET_205;
    wire __A16_NET_206;
    wire __A16_NET_207;
    wire __A16_NET_208;
    wire __A16_NET_209;
    wire __A16_NET_210;
    wire __A16_NET_211;
    wire __A16_NET_212;
    wire __A16_NET_213;
    wire __A16_NET_214;
    wire __A16_NET_215;
    wire __A16_NET_216;
    wire __A16_NET_217;
    wire __A16_NET_218;
    wire __A16_NET_219;
    wire __A16_NET_220;
    wire __A16_NET_221;
    wire __A16_NET_222;
    wire __A16_NET_223;
    wire __A16_NET_224;
    wire __A16_NET_225;
    wire __A16_NET_226;
    wire __A16_NET_227;
    wire __A16_NET_228;
    wire __A16_NET_229;
    wire __A16_NET_230;
    wire __A16_NET_231;
    wire __A16_NET_232;
    wire __A16_NET_233;
    wire __A16_NET_234;
    wire __A16_NET_235;
    wire __A16_NET_236;
    wire __A16_NET_237;
    wire __A16_NET_238;
    wire __A16_NET_239;
    wire __A16_NET_240;
    wire __A16_NET_241;
    wire __A16_NET_242;
    wire __A16_NET_243;
    wire __A16_NET_244;
    wire __A16_NET_245;
    wire __A16_NET_246;
    wire __A16_NET_247;
    wire __A16_NET_248;
    wire __A16_NET_249;
    wire __A16_NET_250;
    wire __A16_NET_251;
    wire __A16_NET_252;
    wire __A16_NET_253;
    wire __A16_NET_254;
    wire __A16_NET_255;
    wire __A16_NET_256;
    wire __A16_NET_257;
    wire __A16_NET_258;
    wire __A16_NET_259;
    wire __A16_NET_260;
    wire __A16_NET_261;
    wire __A16_NET_262;
    wire __A16_NET_263;
    wire __A16_NET_264;
    wire __A16_NET_265;
    wire __A16_NET_266;
    wire __A16_NET_267;
    wire __A16_NET_268;
    wire __A16_NET_269;
    wire __A16_NET_270;
    wire __A16_NET_271;
    wire __A16_NET_272;
    wire __A16_NET_273;

    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16001(__A16_NET_110, CHWL01_n, __A16_1__WCH05_n, __A16_NET_111, __A16_NET_110, __A16_NET_109, GND, __A16_NET_111, __A16_1__CCH05, __A16_NET_109, __A16_NET_111, __A16_1__RCH05_n, __A16_NET_115, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16002(__A16_NET_111, __A16_1__RCpXpP, __A16_NET_112, __A16_1__RCpZpR, __A16_NET_101, __A16_1__RCmXmP, GND, __A16_1__RCmZmR, __A16_NET_106, __A16_1__RCmXpP, __A16_NET_125, __A16_1__RCmZpR, __A16_NET_117, VCC, SIM_RST, SIM_CLK);
    U74HC27 U16003(__A16_NET_104, __A16_NET_115, __A16_NET_121, __A16_NET_105, CH3202, __A16_NET_188, GND, __A16_NET_185, __A16_NET_116, __A16_NET_124, CH3203, __A16_NET_187, CH3201, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U16004(__A16_NET_187, CHOR01_n, __A16_NET_188, CHOR02_n, __A16_NET_185, CHOR03_n, GND, CHOR04_n, __A16_NET_186, CHOR05_n, __A16_NET_191, CHOR06_n, __A16_NET_192, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16005(__A16_NET_114, CHWL01_n, __A16_1__WCH06_n, __A16_NET_112, __A16_NET_114, __A16_NET_113, GND, __A16_NET_112, __A16_1__CCH06, __A16_NET_113, __A16_NET_112, __A16_1__RCH06_n, __A16_NET_104, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16006(__A16_NET_103, CHWL02_n, __A16_1__WCH05_n, __A16_NET_101, __A16_NET_103, __A16_NET_102, GND, __A16_NET_101, __A16_1__CCH05, __A16_NET_102, __A16_NET_101, __A16_1__RCH05_n, __A16_NET_105, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16007(__A16_NET_108, CHWL02_n, __A16_1__WCH06_n, __A16_NET_106, __A16_NET_108, __A16_NET_107, GND, __A16_NET_106, __A16_1__CCH06, __A16_NET_107, __A16_NET_106, __A16_1__RCH06_n, __A16_NET_121, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16008(__A16_NET_127, CHWL03_n, __A16_1__WCH05_n, __A16_NET_125, __A16_NET_127, __A16_NET_126, GND, __A16_NET_125, __A16_1__CCH05, __A16_NET_126, __A16_NET_125, __A16_1__RCH05_n, __A16_NET_124, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16009(__A16_NET_123, CHWL03_n, __A16_1__WCH06_n, __A16_NET_117, __A16_NET_123, __A16_NET_122, GND, __A16_NET_117, __A16_1__CCH06, __A16_NET_122, __A16_NET_117, __A16_1__RCH06_n, __A16_NET_116, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16010(__A16_NET_120, CHWL04_n, __A16_1__WCH05_n, __A16_NET_119, __A16_NET_120, __A16_NET_118, GND, __A16_NET_119, __A16_1__CCH05, __A16_NET_118, __A16_NET_119, __A16_1__RCH05_n, __A16_NET_183, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16011(__A16_NET_119, __A16_1__RCpXmP, __A16_NET_161, __A16_1__RCpZmR, __A16_NET_155, __A16_1__RCpXpY, GND, __A16_1__RCpYpR, __A16_NET_151, __A16_1__RCmXmY, __A16_NET_179, __A16_1__RCmYmR, __A16_NET_184, VCC, SIM_RST, SIM_CLK);
    U74HC27 U16012(__A16_NET_168, __A16_NET_183, __A16_NET_156, __A16_NET_154, CH3205, __A16_NET_191, GND, __A16_NET_192, __A16_NET_182, __A16_NET_178, CH3206, __A16_NET_186, CH3204, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16013(__A16_NET_163, CHWL04_n, __A16_1__WCH06_n, __A16_NET_161, __A16_NET_163, __A16_NET_162, GND, __A16_NET_161, __A16_1__CCH06, __A16_NET_162, __A16_NET_161, __A16_1__RCH06_n, __A16_NET_168, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16014(__A16_NET_165, CHWL05_n, __A16_1__WCH05_n, __A16_NET_155, __A16_NET_165, __A16_NET_164, GND, __A16_NET_155, __A16_1__CCH05, __A16_NET_164, __A16_NET_155, __A16_1__RCH05_n, __A16_NET_154, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16015(__A16_NET_153, CHWL05_n, __A16_1__WCH06_n, __A16_NET_151, __A16_NET_153, __A16_NET_152, GND, __A16_NET_151, __A16_1__CCH06, __A16_NET_152, __A16_NET_151, __A16_1__RCH06_n, __A16_NET_156, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16016(__A16_NET_181, CHWL06_n, __A16_1__WCH05_n, __A16_NET_179, __A16_NET_181, __A16_NET_180, GND, __A16_NET_179, __A16_1__CCH05, __A16_NET_180, __A16_NET_179, __A16_1__RCH05_n, __A16_NET_178, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16017(__A16_NET_177, CHWL06_n, __A16_1__WCH06_n, __A16_NET_184, __A16_NET_177, __A16_NET_176, GND, __A16_NET_184, __A16_1__CCH06, __A16_NET_176, __A16_NET_184, __A16_1__RCH06_n, __A16_NET_182, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16018(__A16_NET_170, CHWL07_n, __A16_1__WCH05_n, __A16_NET_171, __A16_NET_170, __A16_NET_169, GND, __A16_NET_171, __A16_1__CCH05, __A16_NET_169, __A16_NET_171, __A16_1__RCH05_n, __A16_NET_175, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16019(__A16_NET_171, __A16_1__RCmXpY, __A16_NET_172, __A16_1__RCmYpR, __A16_NET_149, __A16_1__RCpXmY, GND, __A16_1__RCpYmR, __A16_NET_145, __A16_1__WCH05_n, __A16_NET_130, __A16_1__WCH06_n, __A16_NET_132, VCC, SIM_RST, SIM_CLK);
    U74HC27 U16020(__A16_NET_144, __A16_NET_175, __A16_NET_142, __A16_NET_148, CH3208, __A16_NET_190, GND, __A16_NET_130, WCHG_n, XT0_n, XB5_n, __A16_NET_189, CH3207, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U16021(__A16_NET_189, CHOR07_n, __A16_NET_190, CHOR08_n, __A16_NET_262, CHOR01_n, GND, CHOR02_n, __A16_NET_259, CHOR03_n, __A16_NET_258, CHOR04_n, __A16_NET_260, VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16022(__A16_NET_174, CHWL07_n, __A16_1__WCH06_n, __A16_NET_172, __A16_NET_174, __A16_NET_173, GND, __A16_NET_172, __A16_1__CCH06, __A16_NET_173, __A16_NET_172, __A16_1__RCH06_n, __A16_NET_144, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16023(__A16_NET_143, CHWL08_n, __A16_1__WCH05_n, __A16_NET_149, __A16_NET_143, __A16_NET_150, GND, __A16_NET_149, __A16_1__CCH05, __A16_NET_150, __A16_NET_149, __A16_1__RCH05_n, __A16_NET_148, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16024(__A16_NET_147, CHWL08_n, __A16_1__WCH06_n, __A16_NET_145, __A16_NET_147, __A16_NET_146, GND, __A16_NET_145, __A16_1__CCH06, __A16_NET_146, __A16_NET_145, __A16_1__RCH06_n, __A16_NET_142, VCC, SIM_RST, SIM_CLK);
    U74HC27 U16025(WCHG_n, XT0_n, CCHG_n, XT0_n, XB5_n, __A16_NET_131, GND, __A16_NET_138, CCHG_n, XT0_n, XB6_n, __A16_NET_132, XB6_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16026(__A16_NET_128, __A16_1__CCH05, __A16_NET_129, __A16_1__RCH05_n, __A16_NET_136, __A16_1__RCH06_n, GND, __A16_1__CCH06, __A16_NET_137, __A16_1__TVCNAB, __A16_NET_139, __A16_1__OT1207, __A16_NET_134, VCC, SIM_RST, SIM_CLK);
    U74HC02 U16027(__A16_NET_128, __A16_NET_131, GOJAM, __A16_NET_129, XT0_n, XB5_n, GND, XT0_n, XB6_n, __A16_NET_136, __A16_NET_138, GOJAM, __A16_NET_137, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16028(__A16_NET_141, CHWL08_n, WCH12_n, __A16_NET_139, __A16_NET_141, __A16_NET_140, GND, __A16_NET_139, CCH12, __A16_NET_140, RCH12_n, __A16_NET_139, CH1208, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16029(__A16_NET_135, WCH12_n, CHWL07_n, __A16_NET_134, __A16_NET_135, __A16_NET_133, GND, __A16_NET_134, CCH12, __A16_NET_133, RCH12_n, __A16_NET_134, __A16_1__CH1207, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16030(__A16_NET_133, __A16_1__OT1207_n, __A16_NET_266, __A16_2__ZOPCDU, __A16_NET_265, __A16_2__ZOPCDU, GND, __A16_2__ENEROP, __A16_NET_225, __A16_2__COMACT, __A16_NET_228, __A16_2__STARON, __A16_NET_217, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16031(__A16_NET_268, CHWL01_n, WCH12_n, __A16_NET_266, __A16_NET_268, __A16_NET_267, GND, __A16_NET_266, CCH12, __A16_NET_267, __A16_NET_266, RCH12_n, __A16_NET_264, VCC, SIM_RST, SIM_CLK);
    U74HC27 U16032(__A16_NET_264, __A16_NET_263, __A16_NET_227, __A16_NET_226, CH1502, __A16_NET_259, GND, __A16_NET_258, __A16_NET_236, __A16_NET_235, CH1503, __A16_NET_262, CH1501, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16033(__A16_NET_269, CHWL01_n, WCH11_n, __A16_NET_265, __A16_NET_269, __A16_NET_261, GND, __A16_NET_265, CCH11, __A16_NET_261, __A16_NET_265, RCH11_n, __A16_NET_263, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16034(__A16_NET_270, CHWL02_n, WCH12_n, __A16_NET_225, __A16_NET_270, __A16_NET_271, GND, __A16_NET_225, CCH12, __A16_NET_271, __A16_NET_225, RCH12_n, __A16_NET_227, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16035(__A16_NET_224, CHWL02_n, WCH11_n, __A16_NET_228, __A16_NET_224, __A16_NET_223, GND, __A16_NET_228, CCH11, __A16_NET_223, __A16_NET_228, RCH11_n, __A16_NET_226, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16036(__A16_NET_219, CHWL03_n, WCH12_n, __A16_NET_217, __A16_NET_219, __A16_NET_218, GND, __A16_NET_217, CCH12, __A16_NET_218, __A16_NET_217, RCH12_n, __A16_NET_236, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16037(__A16_NET_222, CHWL03_n, WCH11_n, __A16_NET_220, __A16_NET_222, __A16_NET_221, GND, __A16_NET_220, CCH11, __A16_NET_221, __A16_NET_220, RCH11_n, __A16_NET_235, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16038(__A16_NET_220, __A16_2__UPLACT, __A16_NET_240, __A16_2__COARSE, __A16_NET_237, TMPOUT, GND, __A16_2__ZIMCDU, __A16_NET_231, __A16_2__ENERIM, __A16_NET_196, __A16_2__S4BTAK, __A16_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16039(__A16_NET_234, CHWL04_n, WCH12_n, __A16_NET_240, __A16_NET_234, __A16_NET_241, GND, __A16_NET_240, CCH12, __A16_NET_241, __A16_NET_240, RCH12_n, __A16_NET_230, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16040(__A16_NET_239, CHWL04_n, WCH11_n, __A16_NET_237, __A16_NET_239, __A16_NET_238, GND, __A16_NET_237, CCH11, __A16_NET_238, __A16_NET_237, RCH11_n, __A16_NET_229, VCC, SIM_RST, SIM_CLK);
    U74HC27 U16041(__A16_NET_230, __A16_NET_229, __A16_NET_199, __A16_NET_205, CH0705, __A16_NET_273, GND, __A16_NET_272, __A16_NET_198, __A16_NET_197, CH0706, __A16_NET_260, CH1504, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16042(__A16_NET_233, CHWL05_n, WCH12_n, __A16_NET_231, __A16_NET_233, __A16_NET_232, GND, __A16_NET_231, CCH12, __A16_NET_232, __A16_NET_231, RCH12_n, __A16_NET_199, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16043(__A16_NET_202, CHWL05_n, WCH11_n, __A16_NET_200, __A16_NET_202, __A16_NET_201, GND, __A16_NET_200, CCH11, __A16_NET_201, __A16_NET_200, RCH11_n, __A16_NET_205, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U16044(__A16_NET_273, CHOR05_n, __A16_NET_272, CHOR06_n, __A16_NET_257, CHOR07_n, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16045(__A16_NET_204, CHWL06_n, WCH12_n, __A16_NET_196, __A16_NET_204, __A16_NET_203, GND, __A16_NET_196, CCH12, __A16_NET_203, __A16_NET_196, RCH12_n, __A16_NET_198, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16046(__A16_NET_195, CHWL06_n, WCH11_n, __A16_NET_193, __A16_NET_195, __A16_NET_194, GND, __A16_NET_193, CCH11, __A16_NET_194, __A16_NET_193, RCH11_n, __A16_NET_197, VCC, SIM_RST, SIM_CLK);
    U74HC02 U16047(__A16_2__KYRLS, __A16_NET_200, FLASH, __A16_2__VNFLSH, __A16_NET_193, FLASH_n, GND, __A16_NET_256, FLASH, __A16_2__OPEROR, __A16_NET_253, GOJAM, __A16_NET_254, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16048(__A16_NET_213, CHWL09_n, WCH12_n, __A16_NET_212, __A16_NET_213, __A16_NET_211, GND, __A16_NET_212, CCH12, __A16_NET_211, __A16_NET_212, RCH12_n, CH1209, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16049(__A16_NET_216, CHWL10_n, WCH12_n, __A16_NET_215, __A16_NET_216, __A16_NET_214, GND, __A16_NET_215, CCH12, __A16_NET_214, __A16_NET_215, RCH12_n, CH1210, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16050(__A16_NET_215, __A16_2__ZEROPT, __A16_NET_207, __A16_2__DISDAC, __A16_NET_247, __A16_2__MROLGT, GND, __A16_2__S4BSEQ, __A16_NET_249, __A16_2__S4BOFF, __A16_NET_242, WCH12_n, __A16_NET_245, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16051(__A16_NET_208, CHWL11_n, WCH12_n, __A16_NET_207, __A16_NET_208, __A16_NET_206, GND, __A16_NET_207, CCH12, __A16_NET_206, __A16_NET_207, RCH12_n, CH1211, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16052(__A16_NET_210, CHWL07_n, WCH11_n, __A16_NET_256, __A16_NET_210, __A16_NET_209, GND, __A16_NET_256, CCH11, __A16_NET_209, __A16_NET_256, RCH11_n, __A16_NET_255, VCC, SIM_RST, SIM_CLK);
    U74HC27 U16053(__A16_1__CH1207, __A16_NET_255, WCHG_n, XB2_n, XT1_n, __A16_NET_245, GND, __A16_NET_253, CCHG_n, XB2_n, XT1_n, __A16_NET_257, CH0707, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16054(__A16_NET_248, CHWL12_n, WCH12_n, __A16_NET_247, __A16_NET_248, __A16_NET_246, GND, __A16_NET_247, CCH12, __A16_NET_246, __A16_NET_247, RCH12_n, CH1212, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16055(__A16_NET_251, CHWL13_n, WCH12_n, __A16_NET_249, __A16_NET_251, __A16_NET_250, GND, __A16_NET_249, CCH12, __A16_NET_250, __A16_NET_249, RCH12_n, CH1213, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16056(__A16_NET_244, CHWL14_n, WCH12_n, __A16_NET_242, __A16_NET_244, __A16_NET_243, GND, __A16_NET_242, CCH12, __A16_NET_243, __A16_NET_242, RCH12_n, CH1214, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16057(__A16_NET_254, CCH12, __A16_NET_252, RCH12_n,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U16058(__A16_NET_252, XT1_n, XB2_n,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
endmodule