`include "components/agc_parts.v"

module stage_branch(VCC, GND, SIM_RST, GOJAM, PHS2_n, PHS3_n, PHS4, PHS4_n, ST1, ST2, T01, T03, T12_n, SQEXT_n, SQ1_n, QC0_n, WL16_n, WL15_n, WL14_n, WL13_n, WL12_n, WL11_n, WL10_n, WL09_n, WL08_n, WL07_n, WL06_n, WL05_n, WL04_n, WL03_n, WL02_n, WL01_n, SUMA16_n, SUMB16_n, DVST, DVST_n, RSTSTG, TOV_n, OVF_n, UNF_n, TSGU_n, TSGN_n, TSGN2, TMZ_n, TPZG_n, GEQZRO_n, TL15, L15_n, TRSM_n, XT1_n, NDR100_n, XB7_n, INKL, STRTFC, ST0_n, ST1_n, STD2, ST3_n, ST4, MTCSAI);
    input wire SIM_RST;
    input wire DVST;
    input wire DVST_n;
    input wire GEQZRO_n;
    input wire GND;
    input wire GOJAM;
    input wire INKL;
    input wire L15_n;
    input wire MTCSAI;
    input wire NDR100_n;
    wire NET_100;
    wire NET_101;
    wire NET_102;
    wire NET_103;
    wire NET_104;
    wire NET_105;
    wire NET_106;
    wire NET_107;
    wire NET_108;
    wire NET_109;
    wire NET_110;
    wire NET_111;
    wire NET_112;
    wire NET_113;
    wire NET_114;
    wire NET_115;
    wire NET_116;
    wire NET_117;
    wire NET_118;
    wire NET_121;
    wire NET_122;
    wire NET_123;
    wire NET_124;
    wire NET_125;
    wire NET_126;
    wire NET_128;
    wire NET_129;
    wire NET_131;
    wire NET_133;
    wire NET_134;
    wire NET_136;
    wire NET_137;
    wire NET_138;
    wire NET_139;
    wire NET_140;
    wire NET_141;
    wire NET_142;
    wire NET_143;
    wire NET_144;
    wire NET_145;
    wire NET_146;
    wire NET_147;
    wire NET_148;
    wire NET_149;
    wire NET_150;
    wire NET_151;
    wire NET_152;
    wire NET_153;
    wire NET_154;
    wire NET_155;
    wire NET_156;
    wire NET_157;
    wire NET_158;
    wire NET_159;
    wire NET_160;
    wire NET_161;
    wire NET_162;
    wire NET_163;
    wire NET_164;
    wire NET_165;
    wire NET_166;
    wire NET_169;
    wire NET_170;
    wire NET_171;
    wire NET_172;
    wire NET_173;
    wire NET_174;
    wire NET_90;
    wire NET_91;
    wire NET_92;
    wire NET_93;
    wire NET_94;
    wire NET_95;
    wire NET_96;
    wire NET_97;
    wire NET_98;
    wire NET_99;
    input wire OVF_n;
    input wire PHS2_n;
    input wire PHS3_n;
    input wire PHS4;
    input wire PHS4_n;
    input wire QC0_n;
    input wire RSTSTG;
    input wire SQ1_n;
    input wire SQEXT_n;
    output wire ST0_n;
    input wire ST1;
    output wire ST1_n;
    input wire ST2;
    output wire ST3_n;
    input wire ST4;
    wire ST4_n;
    output wire STD2;
    input wire STRTFC;
    input wire SUMA16_n;
    input wire SUMB16_n;
    input wire T01;
    input wire T03;
    input wire T12_n;
    input wire TL15;
    input wire TMZ_n;
    input wire TOV_n;
    input wire TPZG_n;
    input wire TRSM_n;
    input wire TSGN2;
    input wire TSGN_n;
    input wire TSGU_n;
    input wire UNF_n;
    input wire VCC;
    input wire WL01_n;
    input wire WL02_n;
    input wire WL03_n;
    input wire WL04_n;
    input wire WL05_n;
    input wire WL06_n;
    input wire WL07_n;
    input wire WL08_n;
    input wire WL09_n;
    input wire WL10_n;
    input wire WL11_n;
    input wire WL12_n;
    input wire WL13_n;
    input wire WL14_n;
    input wire WL15_n;
    input wire WL16_n;
    input wire XB7_n;
    input wire XT1_n;
    wire __A04_1__BR1;
    wire __A04_1__BR1_n;
    wire __A04_1__BR2;
    wire __A04_1__BR2_n;
    wire __A04_1__DIVSTG;
    wire __A04_1__DIV_n;
    wire __A04_1__DV0;
    wire __A04_1__DV0_n;
    wire __A04_1__DV1;
    wire __A04_1__DV1376;
    wire __A04_1__DV1736_n;
    wire __A04_1__DV1_n;
    wire __A04_1__DV376;
    wire __A04_1__DV3764;
    wire __A04_1__DV376_n;
    wire __A04_1__DV4;
    wire __A04_1__MBR1;
    wire __A04_1__MBR2;
    wire __A04_1__MST1;
    wire __A04_1__MST2;
    wire __A04_1__MST3;
    wire __A04_1__SGUM;
    wire __A04_1__ST1376_n;
    wire __A04_1__ST376;
    wire __A04_1__ST376_n;
    wire __A04_1__STG1;
    wire __A04_1__STG2;
    wire __A04_1__STG3;
    wire __A04_1__T12USE_n;

    pullup R2007(NET_118);
    pullup R3004(NET_122);
    pullup R3005(NET_123);
    pullup R4001(NET_156);
    pullup R4002(NET_147);
    pullup R4003(__A04_1__SGUM);
    pullup R4006(NET_129);
    U74HC02 #(0, 0, 0, 1) U4001(__A04_1__T12USE_n, DVST, NET_149, __A04_1__DIVSTG, __A04_1__T12USE_n, T03, GND, NET_150, NET_148, NET_170, GOJAM, MTCSAI, NET_153, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U4002(T03, __A04_1__T12USE_n, __A04_1__T12USE_n, RSTSTG, GOJAM, NET_149, GND, NET_148, PHS3_n, NET_149, T12_n, NET_150, PHS3_n, VCC, SIM_RST);
    U74LVC07 U4003(NET_153, NET_156, NET_155, NET_156, NET_139, NET_147, GND, NET_147, NET_138, __A04_1__SGUM, NET_107, __A04_1__SGUM, NET_106, VCC, SIM_RST);
    U74HC27 #(1, 1, 0) U4004(ST1, NET_151, __A04_1__STG1, __A04_1__STG3, __A04_1__STG2, NET_136, GND, NET_160, __A04_1__STG2, __A04_1__STG3, NET_144, NET_155, NET_154, VCC, SIM_RST);
    U74HC02 U4005(NET_154, NET_156, T01, NET_151, DVST_n, NET_152, GND, NET_170, NET_156, NET_141, NET_154, NET_170, NET_142, VCC, SIM_RST);
    U74HC02 #(1, 0, 1, 0) U4006(NET_144, NET_141, __A04_1__STG1, __A04_1__STG1, NET_144, NET_142, GND, ST2, NET_140, NET_139, DVST_n, NET_144, NET_143, VCC, SIM_RST);
    wire U4007_12_NC;
    wire U4007_13_NC;
    U74HC04 U4007(NET_144, __A04_1__MST1, NET_164, __A04_1__MST2, NET_152, __A04_1__MST3, GND, __A04_1__MBR1, NET_122, __A04_1__MBR2, NET_118, U4007_12_NC, U4007_13_NC, VCC, SIM_RST);
    U74HC04 #(0, 1, 1, 1, 0, 0) U4008(NET_136, ST0_n, NET_160, ST1_n, NET_163, ST3_n, GND, ST4_n, NET_161, __A04_1__ST376_n, __A04_1__ST376, __A04_1__DV1736_n, __A04_1__DV1376, VCC, SIM_RST);
    U74HC27 #(1, 0, 0) U4009(NET_143, MTCSAI, NET_147, GOJAM, T01, NET_137, GND, NET_163, __A04_1__STG3, NET_164, NET_144, NET_138, NET_137, VCC, SIM_RST);
    U74HC4002 U4010(NET_140, TRSM_n, XT1_n, XB7_n, NDR100_n, NET_146, GND, NET_145, NET_174, STRTFC, T01, RSTSTG, NET_165, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U4011(NET_169, NET_170, NET_147, NET_171, NET_137, NET_170, GND, NET_169, __A04_1__STG2, NET_164, NET_164, NET_171, __A04_1__STG2, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U4012(NET_166, DVST_n, NET_164, NET_174, NET_166, NET_165, GND, NET_170, NET_174, NET_172, NET_165, NET_170, NET_173, VCC, SIM_RST);
    U74HC02 #(1, 0, 0, 0) U4013(NET_152, NET_172, __A04_1__STG3, __A04_1__STG3, NET_152, NET_173, GND, __A04_1__STG1, __A04_1__STG3, NET_157, NET_164, NET_157, __A04_1__ST376, VCC, SIM_RST);
    wire U4014_9_NC;
    wire U4014_10_NC;
    wire U4014_11_NC;
    wire U4014_12_NC;
    wire U4014_13_NC;
    U74HC4002 U4014(STD2, INKL, __A04_1__STG1, __A04_1__STG3, NET_164, NET_158, GND, NET_159, U4014_9_NC, U4014_10_NC, U4014_11_NC, U4014_12_NC, U4014_13_NC, VCC, SIM_RST);
    U74HC27 U4015(NET_152, __A04_1__STG1, QC0_n, SQEXT_n, SQ1_n, NET_105, GND, NET_107, SUMB16_n, SUMA16_n, TSGU_n, NET_161, __A04_1__STG2, VCC, SIM_RST);
    U74HC02 U4016(NET_162, NET_161, __A04_1__ST376, __A04_1__DV3764, __A04_1__DIV_n, NET_162, GND, NET_160, __A04_1__ST376, __A04_1__ST1376_n, __A04_1__DIV_n, __A04_1__ST1376_n, __A04_1__DV1376, VCC, SIM_RST);
    U74HC04 U4017(NET_105, __A04_1__DIV_n, __A04_1__DV0, __A04_1__DV0_n, __A04_1__DV1, __A04_1__DV1_n, GND, __A04_1__DV376_n, __A04_1__DV376, NET_94, TL15, __A04_1__BR1, NET_122, VCC, SIM_RST);
    U74HC02 U4018(__A04_1__DV0, __A04_1__DIV_n, ST0_n, __A04_1__DV1, __A04_1__DIV_n, ST1_n, GND, __A04_1__DIV_n, ST4_n, __A04_1__DV4, __A04_1__DIV_n, __A04_1__ST376_n, __A04_1__DV376, VCC, SIM_RST);
    U74HC02 U4019(NET_93, SUMA16_n, SUMB16_n, NET_106, PHS4, PHS3_n, GND, UNF_n, TOV_n, NET_101, L15_n, NET_94, NET_104, VCC, SIM_RST);
    U74HC27 #(0, 0, 1) U4020(PHS4_n, WL16_n, NET_104, NET_103, NET_123, NET_102, GND, NET_97, NET_122, NET_98, NET_90, NET_103, TSGN_n, VCC, SIM_RST);
    U74HC02 U4021(NET_98, TSGN_n, PHS3_n, NET_90, NET_94, PHS3_n, GND, TOV_n, PHS2_n, NET_96, __A04_1__SGUM, NET_101, NET_100, VCC, SIM_RST);
    U74HC4002 U4022(NET_99, NET_93, PHS3_n, TSGU_n, PHS4, NET_92, GND, NET_91, WL16_n, WL15_n, WL14_n, WL13_n, NET_131, VCC, SIM_RST);
    U74LVC07 U4023(NET_100, NET_122, NET_102, NET_122, NET_97, NET_123, GND, NET_123, NET_95, NET_129, NET_131, NET_129, NET_128, VCC, SIM_RST);
    U74HC02 #(1, 0, 0, 0) U4024(NET_95, NET_96, NET_99, NET_115, TOV_n, OVF_n, GND, NET_121, PHS3_n, NET_117, TMZ_n, PHS4_n, NET_113, VCC, SIM_RST);
    wire U4025_10_NC;
    wire U4025_11_NC;
    wire U4025_12_NC;
    wire U4025_13_NC;
    U74HC04 U4025(NET_123, __A04_1__BR1_n, TSGN2, NET_121, NET_118, __A04_1__BR2, GND, __A04_1__BR2_n, NET_110, U4025_10_NC, U4025_11_NC, U4025_12_NC, U4025_13_NC, VCC, SIM_RST);
    U74HC27 U4026(GEQZRO_n, PHS4_n, WL16_n, PHS4_n, NET_121, NET_111, GND, NET_112, NET_111, NET_129, NET_110, NET_108, TPZG_n, VCC, SIM_RST);
    U74HC4002 U4027(NET_128, WL12_n, WL11_n, WL10_n, WL09_n, NET_134, GND, NET_133, WL08_n, WL07_n, WL06_n, WL05_n, NET_126, VCC, SIM_RST);
    U74HC4002 #(0, 1) U4028(NET_114, WL04_n, WL03_n, WL02_n, WL01_n, NET_125, GND, NET_124, NET_118, NET_117, NET_116, NET_96, NET_110, VCC, SIM_RST);
    wire U4029_12_NC;
    wire U4029_13_NC;
    U74LVC07 U4029(NET_126, NET_129, NET_114, NET_129, NET_113, NET_129, GND, NET_118, NET_109, NET_118, NET_112, U4029_12_NC, U4029_13_NC, VCC, SIM_RST);
    wire U4030_8_NC;
    wire U4030_9_NC;
    wire U4030_10_NC;
    wire U4030_11_NC;
    wire U4030_12_NC;
    wire U4030_13_NC;
    U74HC02 U4030(NET_116, TMZ_n, PHS3_n, NET_109, NET_108, NET_115, GND, U4030_8_NC, U4030_9_NC, U4030_10_NC, U4030_11_NC, U4030_12_NC, U4030_13_NC, VCC, SIM_RST);
endmodule