`timescale 1ns/1ps

module crosspoint_ii(VCC, GND, SIM_RST, GOJAM, T01, T01_n, T02, T02_n, T03, T03_n, T04, T04_n, T05, T06, T06_n, T07, T07_n, T08, T08_n, T09, T10, T10_n, T11, T11_n, T12, T12USE_n, PHS4_n, ST2_n, BR1, BR1_n, BR2_n, BR1B2_n, BR12B_n, BR1B2B, BR1B2B_n, INKL, AD0, ADS0, AUG0_n, CCS0, CCS0_n, CDUSTB_n, DAS0, DAS1, DAS1_n, DCA0, DCS0, DIM0_n, DINC, DINC_n, DV1376, DV1376_n, DV376_n, DV4_n, DV4B1B, DXCH0, FETCH1, INCR0, INOTLD, MASK0, MCDU, MINC, MP0T10, MP1, MP1_n, MP3_n, MSU0, NDXX1_n, PCDU, PINC, PRINC, RAND0, RUPT0, RUPT1, SHIFT, STFET1_n, SU0, WAND0, IC6, IC7, IC9, IC11, IC17, B15X, DIVSTG, PTWOX, R6, R15, R1C_n, RADRG, RADRZ, RB1_n, RBSQ, RRPA, STBE, STBF, TL15, L01_n, L02_n, L15_n, MON_n, MONPCH, n8PP4, n1XP10, n2XP3, n2XP5, n2XP7, n2XP8, n3XP2, n3XP6, n3XP7, n4XP11, n5XP4, n5XP12, n5XP15, n5XP21, n5XP28, n6XP5, n6XP8, n7XP4, n7XP9, n7XP19, n8XP6, n9XP1, n9XP5, n10XP1, n10XP8, n11XP2, A2X_n, BXVX, CGMC, CI_n, CLXC, EXT, L2GD_n, MCRO_n, MONEX, MONEX_n, NEAC, PIFL_n, PONEX, R1C, RB_n, RB1, RC_n, RCH_n, RG_n, RU_n, RUS_n, RZ_n, ST1, ST2, TOV_n, TSGU_n, TWOX, WA_n, WB_n, WG_n, WL_n, WQ_n, WS_n, WSC_n, WY_n, WYD_n, WZ_n, ZAP_n, RPTSET, n7XP14);
    input wire SIM_RST;
    inout wire A2X_n;
    input wire AD0;
    input wire ADS0;
    input wire AUG0_n;
    input wire B15X;
    input wire BR1;
    input wire BR12B_n;
    input wire BR1B2B;
    input wire BR1B2B_n;
    input wire BR1B2_n;
    input wire BR1_n;
    input wire BR2_n;
    output wire BXVX;
    input wire CCS0;
    input wire CCS0_n;
    input wire CDUSTB_n;
    output wire CGMC;
    inout wire CI_n;
    output wire CLXC;
    input wire DAS0;
    input wire DAS1;
    input wire DAS1_n;
    input wire DCA0;
    input wire DCS0;
    input wire DIM0_n;
    input wire DINC;
    input wire DINC_n;
    input wire DIVSTG;
    input wire DV1376;
    input wire DV1376_n;
    input wire DV376_n;
    input wire DV4B1B;
    input wire DV4_n;
    input wire DXCH0;
    output wire EXT;
    input wire FETCH1;
    input wire GND;
    input wire GOJAM;
    input wire IC11;
    input wire IC17;
    input wire IC6;
    input wire IC7;
    input wire IC9;
    input wire INCR0;
    input wire INKL;
    input wire INOTLD;
    input wire L01_n;
    input wire L02_n;
    input wire L15_n;
    output wire L2GD_n;
    input wire MASK0;
    input wire MCDU;
    output wire MCRO_n;
    input wire MINC;
    output wire MONEX;
    inout wire MONEX_n;
    input wire MONPCH;
    input wire MON_n;
    input wire MP0T10;
    input wire MP1;
    input wire MP1_n;
    input wire MP3_n;
    input wire MSU0;
    input wire NDXX1_n;
    output wire NEAC;
    wire NET_179;
    wire NET_180;
    wire NET_181;
    wire NET_182;
    wire NET_184;
    wire NET_185;
    wire NET_186;
    wire NET_187;
    wire NET_188;
    wire NET_189;
    wire NET_190;
    wire NET_192;
    wire NET_193;
    wire NET_194;
    wire NET_195;
    wire NET_196;
    wire NET_197;
    wire NET_198;
    wire NET_201;
    wire NET_202;
    wire NET_203;
    wire NET_204;
    wire NET_205;
    wire NET_206;
    wire NET_207;
    wire NET_208;
    wire NET_210;
    wire NET_211;
    wire NET_212;
    wire NET_213;
    wire NET_214;
    wire NET_215;
    wire NET_216;
    wire NET_217;
    wire NET_219;
    wire NET_220;
    wire NET_221;
    wire NET_222;
    wire NET_223;
    wire NET_224;
    wire NET_225;
    wire NET_226;
    wire NET_227;
    wire NET_231;
    wire NET_233;
    wire NET_234;
    wire NET_235;
    wire NET_237;
    wire NET_239;
    wire NET_240;
    wire NET_241;
    wire NET_242;
    wire NET_243;
    wire NET_244;
    wire NET_245;
    wire NET_246;
    wire NET_247;
    wire NET_248;
    wire NET_249;
    wire NET_250;
    wire NET_252;
    wire NET_253;
    wire NET_254;
    wire NET_255;
    wire NET_256;
    wire NET_257;
    wire NET_258;
    wire NET_259;
    wire NET_260;
    wire NET_261;
    wire NET_262;
    wire NET_263;
    wire NET_264;
    wire NET_265;
    wire NET_266;
    wire NET_267;
    wire NET_268;
    wire NET_269;
    wire NET_270;
    wire NET_271;
    wire NET_272;
    wire NET_273;
    wire NET_274;
    wire NET_275;
    wire NET_276;
    wire NET_277;
    wire NET_278;
    wire NET_279;
    wire NET_280;
    wire NET_281;
    wire NET_282;
    wire NET_283;
    wire NET_284;
    wire NET_285;
    wire NET_286;
    wire NET_289;
    wire NET_290;
    wire NET_291;
    wire NET_292;
    wire NET_293;
    wire NET_294;
    wire NET_295;
    wire NET_296;
    wire NET_297;
    wire NET_298;
    wire NET_299;
    wire NET_300;
    wire NET_301;
    wire NET_302;
    wire NET_303;
    wire NET_304;
    wire NET_306;
    wire NET_307;
    wire NET_308;
    wire NET_309;
    wire NET_310;
    wire NET_311;
    wire NET_312;
    wire NET_313;
    wire NET_314;
    wire NET_315;
    wire NET_316;
    wire NET_317;
    wire NET_318;
    wire NET_319;
    wire NET_320;
    wire NET_321;
    wire NET_322;
    wire NET_323;
    wire NET_324;
    wire NET_325;
    wire NET_326;
    wire NET_327;
    wire NET_328;
    wire NET_329;
    wire NET_330;
    wire NET_331;
    wire NET_332;
    wire NET_333;
    wire NET_334;
    wire NET_336;
    wire NET_337;
    wire NET_338;
    wire NET_339;
    wire NET_340;
    input wire PCDU;
    input wire PHS4_n;
    output wire PIFL_n;
    input wire PINC;
    output wire PONEX;
    input wire PRINC;
    input wire PTWOX;
    input wire R15;
    output wire R1C;
    inout wire R1C_n;
    input wire R6;
    input wire RADRG;
    input wire RADRZ;
    input wire RAND0;
    output wire RB1;
    inout wire RB1_n;
    input wire RBSQ;
    inout wire RB_n;
    output wire RCH_n;
    inout wire RC_n;
    inout wire RG_n;
    inout wire RPTSET;
    input wire RRPA;
    input wire RUPT0;
    input wire RUPT1;
    output wire RUS_n;
    inout wire RU_n;
    inout wire RZ_n;
    input wire SHIFT;
    output wire ST1;
    output wire ST2;
    inout wire ST2_n;
    input wire STBE;
    input wire STBF;
    input wire STFET1_n;
    input wire SU0;
    input wire T01;
    input wire T01_n;
    input wire T02;
    input wire T02_n;
    input wire T03;
    input wire T03_n;
    input wire T04;
    input wire T04_n;
    input wire T05;
    input wire T06;
    input wire T06_n;
    input wire T07;
    input wire T07_n;
    input wire T08;
    input wire T08_n;
    input wire T09;
    input wire T10;
    input wire T10_n;
    input wire T11;
    input wire T11_n;
    input wire T12;
    input wire T12USE_n;
    input wire TL15;
    inout wire TOV_n;
    output wire TSGU_n;
    output wire TWOX;
    input wire VCC;
    input wire WAND0;
    inout wire WA_n;
    inout wire WB_n;
    inout wire WG_n;
    inout wire WL_n;
    output wire WQ_n;
    inout wire WSC_n;
    inout wire WS_n;
    inout wire WYD_n;
    inout wire WY_n;
    inout wire WZ_n;
    output wire ZAP_n;
    wire __A06_1__CGMC;
    wire __A06_1__L02A_n;
    wire __A06_1__L15A_n;
    wire __A06_1__RB1F;
    wire __A06_1__ZAP;
    wire __A06_1__ZIP;
    wire __A06_1__ZIPCI;
    wire __A06_2__10XP15;
    wire __A06_2__10XP9;
    wire __A06_2__6XP10;
    wire __A06_2__6XP12;
    wire __A06_2__7XP10;
    wire __A06_2__7XP11;
    wire __A06_2__7XP15;
    wire __A06_2__7XP7;
    wire __A06_2__8XP4;
    wire __A06_2__MOUT;
    wire __A06_2__POUT;
    wire __A06_2__PSEUDO;
    wire __A06_2__RDBANK;
    wire __A06_2__WOVR;
    wire __A06_2__ZOUT;
    input wire n10XP1;
    input wire n10XP8;
    input wire n11XP2;
    input wire n1XP10;
    input wire n2XP3;
    input wire n2XP5;
    input wire n2XP7;
    input wire n2XP8;
    input wire n3XP2;
    input wire n3XP6;
    input wire n3XP7;
    input wire n4XP11;
    input wire n5XP12;
    input wire n5XP15;
    input wire n5XP21;
    input wire n5XP28;
    input wire n5XP4;
    input wire n6XP5;
    input wire n6XP8;
    output wire n7XP14;
    input wire n7XP19;
    input wire n7XP4;
    input wire n7XP9;
    inout wire n8PP4;
    input wire n8XP6;
    input wire n9XP1;
    input wire n9XP5;

    pullup R6001(NET_282);
    pullup R6002(A2X_n);
    pullup R6003(RB_n);
    pullup R6004(WYD_n);
    pullup R6005(NET_267);
    pullup R6006(WL_n);
    pullup R6007(RG_n);
    pullup R6008(WB_n);
    pullup R6009(RU_n);
    pullup R6010(WZ_n);
    pullup R6011(TOV_n);
    pullup R6012(WSC_n);
    pullup R6013(WG_n);
    pullup R6014(NET_217);
    pullup R6015(NET_220);
    pullup R6016(MONEX_n);
    pullup R6017(RB1_n);
    pullup R6018(R1C_n);
    pullup R6019(n8PP4);
    pullup R6020(NET_204);
    pullup R6021(WS_n);
    pullup R6022(NET_206);
    pullup R6023(CI_n);
    pullup R6024(WA_n);
    pullup R6025(NET_241);
    pullup R6026(ST2_n);
    pullup R6027(RZ_n);
    pullup R6028(RC_n);
    U74HC27 U6001(T04, T07, NET_279, NET_280, NET_281, NET_286, GND, NET_298, T01, T03, T05, NET_285, T10, VCC, SIM_RST);
    U74HC02 U6002(NET_279, NET_285, DV376_n, NET_280, T01_n, DV1376_n, GND, T04_n, DV4_n, NET_281, MP1_n, NET_282, NET_283, VCC, SIM_RST);
    U74HC27 #(0, 0, 1) U6003(T07, T09, __A06_1__L15A_n, __A06_1__L02A_n, L01_n, NET_333, GND, NET_339, T05, T08, T11, NET_297, T11, VCC, SIM_RST);
    U74LVC07 U6004(NET_298, NET_282, NET_297, NET_282, NET_296, A2X_n, GND, RB_n, NET_308, WYD_n, NET_311, WY_n, NET_301, VCC, SIM_RST);
    U74HC02 #(1, 0, 1, 0) U6005(NET_307, NET_283, n2XP7, L2GD_n, __A06_1__ZIP, CGMC, GND, CGMC, NET_300, NET_311, NET_299, NET_302, NET_303, VCC, SIM_RST);
    U74HC04 U6006(L01_n, NET_310, __A06_1__L02A_n, NET_332, __A06_1__L15A_n, NET_331, GND, CGMC, NET_286, __A06_1__ZIP, NET_307, NET_336, NET_334, VCC, SIM_RST);
    U74HC27 #(1, 0, 0) U6007(n7XP19, __A06_1__ZIP, CGMC, NET_304, RBSQ, NET_308, GND, NET_309, NET_310, NET_332, NET_331, NET_296, CGMC, VCC, SIM_RST);
    U74HC27 U6008(NET_331, NET_310, NET_307, NET_302, NET_299, NET_321, GND, NET_334, NET_299, NET_302, __A06_1__L02A_n, NET_302, __A06_1__L02A_n, VCC, SIM_RST);
    U74HC02 U6009(NET_300, NET_307, NET_303, NET_306, NET_307, NET_336, GND, NET_339, DV376_n, NET_273, DV1376_n, T02_n, NET_271, VCC, SIM_RST);
    U74HC04 U6010(NET_306, MCRO_n, NET_272, NET_269, NET_278, NET_275, GND, __A06_1__ZAP, ZAP_n, NET_317, NET_339, MONEX, MONEX_n, VCC, SIM_RST);
    U74HC27 U6011(NET_307, NET_336, NET_334, NET_309, NET_307, NET_304, GND, NET_299, NET_332, __A06_1__L15A_n, L01_n, __A06_1__ZIPCI, NET_333, VCC, SIM_RST);
    U74HC02 #(1, 1, 1, 0) U6012(NET_272, NET_273, NET_271, NET_278, NET_277, DIVSTG, GND, T08, T10, NET_265, MP1_n, NET_267, NET_266, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U6013(T06, T09, DV376_n, NET_276, T12USE_n, NET_277, GND, NET_274, T02, T04, T06, NET_276, T12, VCC, SIM_RST);
    U74LVC07 U6014(NET_274, NET_267, NET_265, NET_267, NET_268, WL_n, GND, RG_n, NET_290, WB_n, NET_289, RU_n, NET_293, VCC, SIM_RST);
    U74HC02 #(1, 0, 1, 0) U6015(NET_264, T01, T03, NET_270, NET_264, MP3_n, GND, NET_266, NET_270, ZAP_n, n5XP28, NET_269, TSGU_n, VCC, SIM_RST);
    U74HC02 #(1, 1, 1, 0) U6016(NET_268, NET_269, n5XP12, NET_284, RRPA, n5XP4, GND, n5XP15, n3XP6, WQ_n, n9XP5, n6XP8, NET_338, VCC, SIM_RST);
    U74HC4002 #(0, 1) U6017(NET_290, n5XP4, RADRG, NET_269, n5XP28, NET_291, GND, NET_292, n5XP28, n1XP10, NET_275, n2XP3, NET_289, VCC, SIM_RST);
    U74HC4002 U6018(NET_293, NET_275, __A06_1__ZAP, n5XP12, n6XP5, NET_294, GND, NET_295, PRINC, PINC, MINC, DINC, NET_231, VCC, SIM_RST);
    U74LVC07 U6019(NET_284, WZ_n, NET_340, TOV_n, NET_338, WSC_n, GND, WG_n, NET_337, NET_217, NET_262, NET_217, NET_263, VCC, SIM_RST);
    U74HC27 U6020(n6XP5, n3XP2, BR1_n, PHS4_n, TSGU_n, __A06_1__RB1F, GND, CLXC, TSGU_n, BR1, PHS4_n, NET_340, n9XP5, VCC, SIM_RST);
    U74HC02 #(0, 1, 1, 1) U6021(NET_337, n6XP8, n6XP8, PIFL_n, CGMC, NET_318, GND, PTWOX, MONEX, NET_313, MONEX, B15X, NET_314, VCC, SIM_RST);
    U74HC27 U6022(PIFL_n, NET_317, STBE, n1XP10, STBF, NET_312, GND, NET_262, NET_261, NET_260, INCR0, NET_318, T02, VCC, SIM_RST);
    U74HC04 U6023(NET_313, TWOX, NET_314, BXVX, NET_330, NET_316, GND, NET_327, NET_316, NET_328, NET_327, NET_326, NET_328, VCC, SIM_RST);
    U74HC02 U6024(__A06_1__CGMC, NET_312, NET_330, NET_315, __A06_1__CGMC, NET_324, GND, NET_315, NET_312, NET_330, BR1, AUG0_n, NET_261, VCC, SIM_RST);
    U74HC04 #(0, 0, 0, 0, 1, 0) U6025(NET_326, NET_322, NET_322, NET_323, NET_323, NET_325, GND, NET_324, NET_325, NET_210, NET_221, NET_235, __A06_2__7XP10, VCC, SIM_RST);
    U74HC02 U6026(NET_260, DIM0_n, BR12B_n, NET_263, PINC, NET_257, GND, BR12B_n, DINC_n, NET_257, T06_n, NET_217, __A06_2__6XP10, VCC, SIM_RST);
    U74HC02 U6027(NET_215, MINC, MCDU, NET_222, AUG0_n, BR1_n, GND, DIM0_n, BR1B2B_n, NET_223, BR1B2B_n, DINC_n, NET_219, VCC, SIM_RST);
    U74HC27 U6028(NET_222, NET_223, BR1B2B_n, CDUSTB_n, DINC_n, __A06_2__POUT, GND, __A06_2__MOUT, BR12B_n, CDUSTB_n, DINC_n, NET_216, NET_219, VCC, SIM_RST);
    U74LVC07 U6029(NET_215, NET_220, NET_216, NET_220, NET_210, MONEX_n, GND, WA_n, NET_212, RB1_n, NET_235, R1C_n, NET_225, VCC, SIM_RST);
    U74HC02 U6030(NET_221, T06_n, NET_220, NET_211, PCDU, MCDU, GND, T06_n, NET_211, __A06_2__6XP12, NET_213, T07_n, NET_214, VCC, SIM_RST);
    U74HC27 #(0, 1, 1) U6031(BR2_n, DINC_n, DAS0, DAS1, MSU0, NET_213, GND, NET_212, NET_214, __A06_2__7XP7, NET_205, __A06_2__ZOUT, CDUSTB_n, VCC, SIM_RST);
    U74HC02 U6032(NET_233, DV4_n, BR1B2B, __A06_2__7XP7, T07_n, NET_234, GND, WAND0, INOTLD, NET_237, T07_n, NET_237, n7XP14, VCC, SIM_RST);
    U74HC27 U6033(NET_233, WAND0, DAS1_n, T07_n, BR1B2_n, __A06_2__7XP10, GND, __A06_2__7XP11, DAS1_n, T07_n, BR12B_n, NET_234, RAND0, VCC, SIM_RST);
    U74HC04 U6034(__A06_2__7XP11, NET_225, NET_196, PONEX, ST2_n, ST2, GND, ST1, NET_249, NET_246, __A06_2__PSEUDO, NET_247, __A06_2__RDBANK, VCC, SIM_RST);
    U74HC02 U6035(__A06_2__7XP15, NET_224, T07_n, NET_227, NET_231, T07_n, GND, PRINC, INKL, NET_188, IC9, DXCH0, NET_190, VCC, SIM_RST);
    U74HC27 U6036(PCDU, MCDU, n7XP9, n11XP2, __A06_2__7XP15, RUS_n, GND, NET_226, NET_227, NET_239, NET_205, NET_224, SHIFT, VCC, SIM_RST);
    U74LVC07 U6037(NET_226, RU_n, NET_186, WSC_n, NET_189, WG_n, GND, RB_n, NET_181, n8PP4, NET_182, n8PP4, NET_179, VCC, SIM_RST);
    U74HC27 U6038(NET_188, T07_n, T04_n, MON_n, FETCH1, NET_187, GND, NET_186, __A06_2__WOVR, NET_187, NET_192, __A06_2__WOVR, MONPCH, VCC, SIM_RST);
    U74HC02 U6039(NET_189, __A06_2__WOVR, NET_192, NET_192, T07_n, NET_190, GND, __A06_2__10XP9, NET_192, NET_181, T08_n, n8PP4, __A06_2__8XP4, VCC, SIM_RST);
    U74HC27 U6040(RUPT1, DAS1, IC17, MASK0, IC11, NET_179, GND, NET_180, IC6, IC7, IC9, NET_182, MSU0, VCC, SIM_RST);
    U74LVC07 U6041(NET_180, n8PP4, NET_184, NET_204, NET_185, NET_204, GND, WS_n, NET_203, NET_206, NET_207, NET_206, NET_195, VCC, SIM_RST);
    U74HC27 U6042(T08_n, RUPT0, NET_204, R6, R15, NET_203, GND, NET_195, ADS0, IC11, NET_197, NET_184, DAS0, VCC, SIM_RST);
    U74HC02 U6043(NET_185, MP1, DV1376, NET_208, MP3_n, BR1_n, GND, NET_208, CCS0, NET_207, T11_n, NET_206, NET_205, VCC, SIM_RST);
    U74HC02 U6044(NET_197, DAS1_n, BR2_n, NET_202, __A06_1__ZIPCI, __A06_2__6XP12, GND, CCS0_n, BR1B2B_n, NET_198, T10_n, NDXX1_n, EXT, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U6045(T03_n, DAS1_n, NET_244, NET_239, n2XP5, NET_256, GND, NET_254, IC7, DCS0, SU0, NET_239, ADS0, VCC, SIM_RST);
    U74HC4002 #(1, 0) U6046(NET_196, n8XP6, n7XP4, n10XP8, __A06_2__6XP10, NET_193, GND, NET_194, IC6, DCA0, AD0, NET_198, NET_201, VCC, SIM_RST);
    U74LVC07 U6047(NET_202, CI_n, NET_256, WA_n, NET_253, RC_n, GND, NET_241, NET_254, NET_241, NET_252, ST2_n, NET_255, VCC, SIM_RST);
    U74HC02 U6048(__A06_2__10XP9, T10_n, NET_201, NET_243, IC6, IC7, GND, T10_n, NET_243, NET_244, T10_n, NET_241, NET_240, VCC, SIM_RST);
    U74HC02 U6049(NET_253, NET_240, __A06_2__7XP7, NET_252, NET_242, DV4B1B, GND, CCS0_n, BR12B_n, NET_242, T10_n, MP1_n, __A06_2__10XP15, VCC, SIM_RST);
    U74HC27 U6050(__A06_2__8XP4, __A06_2__10XP15, __A06_2__8XP4, RADRZ, n9XP1, NET_248, GND, NEAC, NET_250, TL15, GOJAM, NET_255, RADRZ, VCC, SIM_RST);
    wire U6051_9_NC;
    wire U6051_10_NC;
    wire U6051_11_NC;
    wire U6051_12_NC;
    wire U6051_13_NC;
    U74HC4002 U6051(NET_249, n2XP8, n10XP1, MP0T10, __A06_2__10XP15, NET_258, GND, NET_259, U6051_9_NC, U6051_10_NC, U6051_11_NC, U6051_12_NC, U6051_13_NC, VCC, SIM_RST);
    wire U6052_10_NC;
    wire U6052_11_NC;
    wire U6052_12_NC;
    wire U6052_13_NC;
    U74LVC07 U6052(NET_248, RZ_n, NET_246, RPTSET, NET_247, RU_n, GND, RC_n, NET_329, U6052_10_NC, U6052_11_NC, U6052_12_NC, U6052_13_NC, VCC, SIM_RST);
    U74HC02 #(1, 0, 0, 0) U6053(NET_250, MP0T10, NEAC, NET_245, RADRZ, __A06_2__PSEUDO, GND, T06_n, STFET1_n, __A06_2__RDBANK, __A06_1__ZIPCI, n3XP7, NET_329, VCC, SIM_RST);
    wire U6054_8_NC;
    wire U6054_9_NC;
    wire U6054_10_NC;
    wire U6054_11_NC;
    U74HC27 #(1, 0, 0) U6054(NET_245, GOJAM, n3XP7, n5XP21, n4XP11, RCH_n, GND, U6054_8_NC, U6054_9_NC, U6054_10_NC, U6054_11_NC, __A06_2__PSEUDO, RADRG, VCC, SIM_RST);
    U74HC04 #(0, 0, 0, 1, 0, 0) U6055(R1C_n, R1C, RB1_n, RB1, L02_n, NET_320, GND, __A06_1__L02A_n, NET_320, NET_319, L15_n, __A06_1__L15A_n, NET_319, VCC, SIM_RST);
    wire U6056_3_NC;
    wire U6056_4_NC;
    wire U6056_5_NC;
    wire U6056_6_NC;
    wire U6056_8_NC;
    wire U6056_9_NC;
    wire U6056_10_NC;
    wire U6056_11_NC;
    wire U6056_12_NC;
    wire U6056_13_NC;
    U74HC04 #(1, 0, 0, 0, 0, 0) U6056(NET_321, NET_301, U6056_3_NC, U6056_4_NC, U6056_5_NC, U6056_6_NC, GND, U6056_8_NC, U6056_9_NC, U6056_10_NC, U6056_11_NC, U6056_12_NC, U6056_13_NC, VCC, SIM_RST);
endmodule