`timescale 1ns/1ps
`default_nettype none

module inout_v(SIM_RST, SIM_CLK, p4VDC, p4VSW, GND, GOJAM, T10_n, F10A, CCH13, CCH33, CCH34, CCH35, RCH13_n, RCH33_n, WCH13_n, WCH34_n, WCH35_n, DKSTRT, DKEND, DKBSNC, DRPRST, PC15_n, CHWL01_n, CHWL02_n, CHWL03_n, CHWL04_n, CHWL05_n, CHWL06_n, CHWL07_n, CHWL08_n, CHWL09_n, CHWL10_n, CHWL11_n, CHWL12_n, CHWL13_n, CHWL14_n, CHWL16_n, DLKPLS, CH1307, CH3312);
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire p4VDC;
    input wire p4VSW;
    input wire GND;
    input wire CCH13;
    input wire CCH33;
    input wire CCH34;
    input wire CCH35;
    output wire CH1307;
    output wire CH3312;
    input wire CHWL01_n;
    input wire CHWL02_n;
    input wire CHWL03_n;
    input wire CHWL04_n;
    input wire CHWL05_n;
    input wire CHWL06_n;
    input wire CHWL07_n;
    input wire CHWL08_n;
    input wire CHWL09_n;
    input wire CHWL10_n;
    input wire CHWL11_n;
    input wire CHWL12_n;
    input wire CHWL13_n;
    input wire CHWL14_n;
    input wire CHWL16_n;
    input wire DKBSNC;
    input wire DKEND;
    input wire DKSTRT;
    output wire DLKPLS;
    input wire DRPRST;
    input wire F10A;
    input wire GOJAM;
    input wire PC15_n;
    input wire RCH13_n;
    input wire RCH33_n;
    input wire T10_n;
    input wire WCH13_n;
    input wire WCH34_n;
    input wire WCH35_n;
    wire __A22_1__16CNT;
    wire __A22_1__1CNT;
    wire __A22_1__32CNT;
    wire __A22_1__ADVCTR;
    wire __A22_1__BSYNC_n;
    wire __A22_1__DATA_n; //FPGA#wand
    wire __A22_1__DKCTR1;
    wire __A22_1__DKCTR1_n;
    wire __A22_1__DKCTR2;
    wire __A22_1__DKCTR2_n;
    wire __A22_1__DKCTR3;
    wire __A22_1__DKCTR3_n;
    wire __A22_1__DKCTR4;
    wire __A22_1__DKCTR4_n;
    wire __A22_1__DKCTR5;
    wire __A22_1__DKCTR5_n;
    wire __A22_1__DKDATA;
    wire __A22_1__DKDATB;
    wire __A22_1__DKDAT_n;
    wire __A22_1__DLKCLR;
    wire __A22_1__DLKRPT;
    wire __A22_1__END;
    wire __A22_1__HIGH0_n;
    wire __A22_1__HIGH1_n;
    wire __A22_1__HIGH2_n;
    wire __A22_1__HIGH3_n;
    wire __A22_1__LOW0_n;
    wire __A22_1__LOW1_n;
    wire __A22_1__LOW2_n;
    wire __A22_1__LOW3_n;
    wire __A22_1__LOW4_n;
    wire __A22_1__LOW5_n;
    wire __A22_1__LOW6_n;
    wire __A22_1__LOW7_n;
    wire __A22_1__ORDRBT;
    wire __A22_1__RDOUT_n;
    wire __A22_1__WDORDR;
    wire __A22_1__WRD1B1;
    wire __A22_1__WRD1BP;
    wire __A22_1__WRD2B2;
    wire __A22_1__WRD2B3;
    wire __A22_NET_101;
    wire __A22_NET_102;
    wire __A22_NET_103;
    wire __A22_NET_104;
    wire __A22_NET_105;
    wire __A22_NET_106;
    wire __A22_NET_108;
    wire __A22_NET_109;
    wire __A22_NET_110;
    wire __A22_NET_112;
    wire __A22_NET_113;
    wire __A22_NET_117;
    wire __A22_NET_118;
    wire __A22_NET_119;
    wire __A22_NET_120;
    wire __A22_NET_121;
    wire __A22_NET_122;
    wire __A22_NET_123;
    wire __A22_NET_124;
    wire __A22_NET_125;
    wire __A22_NET_126;
    wire __A22_NET_128;
    wire __A22_NET_129;
    wire __A22_NET_130;
    wire __A22_NET_131;
    wire __A22_NET_132;
    wire __A22_NET_133;
    wire __A22_NET_134;
    wire __A22_NET_136;
    wire __A22_NET_137;
    wire __A22_NET_138;
    wire __A22_NET_139;
    wire __A22_NET_140;
    wire __A22_NET_141;
    wire __A22_NET_142;
    wire __A22_NET_143;
    wire __A22_NET_144;
    wire __A22_NET_145;
    wire __A22_NET_146;
    wire __A22_NET_147;
    wire __A22_NET_148;
    wire __A22_NET_149;
    wire __A22_NET_150;
    wire __A22_NET_151;
    wire __A22_NET_152;
    wire __A22_NET_153;
    wire __A22_NET_154;
    wire __A22_NET_155;
    wire __A22_NET_156;
    wire __A22_NET_157;
    wire __A22_NET_158;
    wire __A22_NET_159;
    wire __A22_NET_160;
    wire __A22_NET_161;
    wire __A22_NET_162;
    wire __A22_NET_163;
    wire __A22_NET_164;
    wire __A22_NET_165;
    wire __A22_NET_168;
    wire __A22_NET_169;
    wire __A22_NET_170;
    wire __A22_NET_171;
    wire __A22_NET_172;
    wire __A22_NET_173;
    wire __A22_NET_174;
    wire __A22_NET_175;
    wire __A22_NET_176;
    wire __A22_NET_177;
    wire __A22_NET_178;
    wire __A22_NET_181;
    wire __A22_NET_182;
    wire __A22_NET_183;
    wire __A22_NET_184;
    wire __A22_NET_185;
    wire __A22_NET_186;
    wire __A22_NET_187;
    wire __A22_NET_188;
    wire __A22_NET_189;
    wire __A22_NET_190;
    wire __A22_NET_191;
    wire __A22_NET_192;
    wire __A22_NET_193;
    wire __A22_NET_194;
    wire __A22_NET_195;
    wire __A22_NET_196;
    wire __A22_NET_197;
    wire __A22_NET_198;
    wire __A22_NET_199;
    wire __A22_NET_200;
    wire __A22_NET_201;
    wire __A22_NET_202;
    wire __A22_NET_203;
    wire __A22_NET_204;
    wire __A22_NET_205;
    wire __A22_NET_206;
    wire __A22_NET_207;
    wire __A22_NET_208;
    wire __A22_NET_209;
    wire __A22_NET_210;
    wire __A22_NET_211;
    wire __A22_NET_212;
    wire __A22_NET_214;
    wire __A22_NET_215;
    wire __A22_NET_216;
    wire __A22_NET_218;
    wire __A22_NET_219;
    wire __A22_NET_220;
    wire __A22_NET_221;
    wire __A22_NET_222;
    wire __A22_NET_223;
    wire __A22_NET_224;
    wire __A22_NET_225;
    wire __A22_NET_226;
    wire __A22_NET_227;
    wire __A22_NET_228;
    wire __A22_NET_229;
    wire __A22_NET_230;
    wire __A22_NET_231;
    wire __A22_NET_232;
    wire __A22_NET_233;
    wire __A22_NET_234;
    wire __A22_NET_235;
    wire __A22_NET_236;
    wire __A22_NET_237;
    wire __A22_NET_238;
    wire __A22_NET_239;
    wire __A22_NET_240;
    wire __A22_NET_241;
    wire __A22_NET_242;
    wire __A22_NET_243;
    wire __A22_NET_244;
    wire __A22_NET_245;
    wire __A22_NET_246;
    wire __A22_NET_247;
    wire __A22_NET_248;
    wire __A22_NET_249;
    wire __A22_NET_252;
    wire __A22_NET_253;
    wire __A22_NET_254;
    wire __A22_NET_255;
    wire __A22_NET_256;
    wire __A22_NET_257;
    wire __A22_NET_258;
    wire __A22_NET_259;
    wire __A22_NET_260;
    wire __A22_NET_262;
    wire __A22_NET_263;
    wire __A22_NET_264;
    wire __A22_NET_266;
    wire __A22_NET_267;
    wire __A22_NET_268;
    wire __A22_NET_269;
    wire __A22_NET_270;
    wire __A22_NET_271;
    wire __A22_NET_272;
    wire __A22_NET_273;
    wire __A22_NET_274;
    wire __A22_NET_275;
    wire __A22_NET_276;
    wire __A22_NET_277;
    wire __A22_NET_280;
    wire __A22_NET_281;
    wire __A22_NET_282;
    wire __A22_NET_283;
    wire __A22_NET_284;
    wire __A22_NET_285;
    wire __A22_NET_286;
    wire __A22_NET_287;
    wire __A22_NET_288;
    wire __A22_NET_54;
    wire __A22_NET_59;
    wire __A22_NET_60;
    wire __A22_NET_61;
    wire __A22_NET_64;
    wire __A22_NET_66;
    wire __A22_NET_67;
    wire __A22_NET_68;
    wire __A22_NET_69;
    wire __A22_NET_71;
    wire __A22_NET_74;
    wire __A22_NET_75;
    wire __A22_NET_78;
    wire __A22_NET_79;
    wire __A22_NET_80;
    wire __A22_NET_81;
    wire __A22_NET_82;
    wire __A22_NET_83;
    wire __A22_NET_84;
    wire __A22_NET_85;
    wire __A22_NET_86;
    wire __A22_NET_87;
    wire __A22_NET_88;
    wire __A22_NET_89;
    wire __A22_NET_90;
    wire __A22_NET_93;
    wire __A22_NET_95;
    wire __A22_NET_99;

    pullup R22001(__A22_1__DATA_n);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0) U22001(__A22_NET_129, __A22_1__DLKRPT, __A22_NET_128, DLKPLS, T10_n, __A22_NET_129, GND, __A22_NET_134, __A22_NET_125, __A22_1__DLKRPT, __A22_1__DLKRPT, __A22_NET_124, __A22_NET_125, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22002(__A22_NET_129, DRPRST, __A22_NET_134, __A22_1__DLKRPT, __A22_NET_124, __A22_NET_130, GND, __A22_1__ADVCTR, __A22_1__RDOUT_n, __A22_1__WDORDR, __A22_1__BSYNC_n, __A22_NET_128, GOJAM, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0) U22003(DKEND, __A22_NET_134, __A22_NET_134, __A22_1__END, DKSTRT, __A22_NET_133, GND, __A22_1__DLKCLR, __A22_NET_133, __A22_NET_112, __A22_NET_110, __A22_1__DKCTR1_n, __A22_NET_118, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b0) U22004(__A22_NET_124, __A22_1__DLKRPT, __A22_NET_126, __A22_NET_126, __A22_NET_124, F10A, GND, __A22_NET_130, __A22_NET_132, __A22_NET_131, __A22_NET_131, CCH33, __A22_NET_132, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0, 1'b0) U22005(CH3312, RCH33_n, __A22_NET_132, __A22_NET_110, __A22_1__DLKCLR, __A22_1__ADVCTR, GND, __A22_1__DLKCLR, __A22_NET_113, __A22_1__RDOUT_n, __A22_1__RDOUT_n, __A22_1__END, __A22_NET_113, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0, 1'b0) U22006(__A22_1__1CNT, __A22_NET_112, __A22_NET_122, __A22_NET_112, __A22_NET_119, __A22_NET_123, GND, __A22_NET_117, __A22_NET_118, __A22_1__DLKCLR, __A22_NET_123, __A22_NET_122, __A22_NET_123, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1, 1'b0) U22007(__A22_1__1CNT, __A22_NET_118, __A22_NET_122, __A22_NET_119, __A22_NET_123, __A22_NET_117, GND, __A22_NET_122, __A22_NET_117, __A22_NET_118, __A22_NET_147, __A22_NET_120, __A22_NET_121, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U22008(__A22_NET_117, __A22_1__DKCTR1, __A22_NET_147, __A22_1__DKCTR2_n, __A22_NET_148, __A22_1__DKCTR2, GND, __A22_1__DKCTR3_n, __A22_NET_138, __A22_1__DKCTR3, __A22_NET_139, __A22_1__DKCTR4_n, __A22_NET_145, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0, 1'b0) U22009(__A22_NET_121, __A22_NET_119, __A22_NET_120, __A22_NET_119, __A22_NET_151, __A22_NET_149, GND, __A22_NET_148, __A22_NET_147, __A22_1__DLKCLR, __A22_NET_149, __A22_NET_120, __A22_NET_149, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0, 1'b0) U22010(__A22_NET_151, __A22_NET_149, __A22_NET_148, __A22_NET_147, __A22_NET_120, __A22_NET_148, GND, __A22_NET_138, __A22_NET_152, __A22_NET_150, __A22_NET_153, __A22_NET_139, __A22_NET_140, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0, 1'b0) U22011(__A22_NET_150, __A22_NET_151, __A22_NET_152, __A22_NET_151, __A22_NET_140, __A22_NET_153, GND, __A22_NET_139, __A22_NET_138, __A22_1__DLKCLR, __A22_NET_153, __A22_NET_152, __A22_NET_153, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b0, 1'b1, 1'b0) U22012(__A22_NET_138, __A22_NET_152, __A22_NET_139, __A22_NET_136, __A22_NET_145, __A22_NET_137, GND, __A22_NET_144, __A22_NET_146, __A22_NET_141, __A22_NET_137, __A22_NET_146, __A22_NET_145, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0, 1'b0) U22013(__A22_NET_136, __A22_NET_140, __A22_NET_137, __A22_NET_140, __A22_NET_141, __A22_NET_144, GND, __A22_NET_146, __A22_NET_145, __A22_1__DLKCLR, __A22_NET_144, __A22_NET_137, __A22_NET_144, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0) U22014(__A22_NET_146, __A22_1__DKCTR4, __A22_NET_74, __A22_1__DKCTR5_n, __A22_NET_75, __A22_1__DKCTR5, GND, __A22_NET_85, __A22_1__BSYNC_n, __A22_NET_84, __A22_NET_83, __A22_NET_79, __A22_NET_84, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b0) U22015(__A22_1__16CNT, __A22_NET_74, __A22_NET_142, __A22_1__32CNT, __A22_NET_143, __A22_NET_75, GND, __A22_NET_142, __A22_NET_75, __A22_NET_74, __A22_NET_85, __A22_NET_79, __A22_NET_82, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0, 1'b0) U22016(__A22_1__16CNT, __A22_NET_141, __A22_NET_142, __A22_NET_141, __A22_1__32CNT, __A22_NET_143, GND, __A22_NET_75, __A22_NET_74, __A22_1__DLKCLR, __A22_NET_143, __A22_NET_142, __A22_NET_143, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U22017(__A22_NET_78, __A22_NET_82, __A22_NET_83, __A22_NET_83, __A22_NET_85, __A22_NET_78, GND, CHWL07_n, WCH13_n, __A22_NET_80, __A22_NET_81, __A22_NET_80, __A22_NET_64, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b0) U22018(__A22_NET_81, CCH13, __A22_NET_64, CH1307, RCH13_n, __A22_NET_64, GND, __A22_1__DLKCLR, __A22_1__WDORDR, __A22_NET_60, __A22_NET_60, __A22_NET_82, __A22_1__WDORDR, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U22019(__A22_1__ORDRBT, __A22_NET_64, __A22_NET_60, __A22_NET_59, __A22_1__DKCTR5, __A22_1__DKCTR4, GND, __A22_1__DKCTR5, __A22_1__DKCTR4_n, __A22_NET_61, __A22_1__DKCTR4, __A22_1__DKCTR5_n, __A22_NET_69, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U22020(__A22_NET_59, __A22_1__HIGH0_n, __A22_NET_61, __A22_1__HIGH1_n, __A22_NET_69, __A22_1__HIGH2_n, GND, __A22_1__HIGH3_n, __A22_NET_71, __A22_1__LOW0_n, __A22_NET_67, __A22_1__LOW1_n, __A22_NET_66, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U22021(__A22_NET_71, __A22_1__DKCTR4_n, __A22_1__DKCTR5_n, __A22_NET_102, CHWL16_n, WCH34_n, GND, __A22_NET_102, __A22_NET_104, __A22_NET_103, __A22_NET_103, CCH34, __A22_NET_104, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22022(__A22_1__DKCTR1, __A22_1__DKCTR2, __A22_1__DKCTR1_n, __A22_1__DKCTR2, __A22_1__DKCTR3, __A22_NET_66, GND, __A22_NET_68, __A22_1__DKCTR1, __A22_1__DKCTR2_n, __A22_1__DKCTR3, __A22_NET_67, __A22_1__DKCTR3, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U22023(__A22_NET_68, __A22_1__LOW2_n, __A22_NET_101, __A22_1__LOW3_n, __A22_NET_95, __A22_1__LOW4_n, GND, __A22_1__LOW5_n, __A22_NET_99, __A22_1__LOW6_n, __A22_NET_108, __A22_1__LOW7_n, __A22_NET_109, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22024(__A22_1__DKCTR1_n, __A22_1__DKCTR2_n, __A22_1__DKCTR1, __A22_1__DKCTR2, __A22_1__DKCTR3_n, __A22_NET_95, GND, __A22_NET_99, __A22_1__DKCTR1_n, __A22_1__DKCTR2, __A22_1__DKCTR3_n, __A22_NET_101, __A22_1__DKCTR3, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22025(__A22_1__DKCTR1, __A22_1__DKCTR2_n, __A22_1__DKCTR1_n, __A22_1__DKCTR2_n, __A22_1__DKCTR3_n, __A22_NET_109, GND, __A22_NET_88, __A22_1__LOW0_n, __A22_NET_103, __A22_1__HIGH0_n, __A22_NET_108, __A22_1__DKCTR3_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U22026(__A22_NET_105, WCH34_n, CHWL14_n, __A22_NET_90, __A22_NET_105, __A22_NET_106, GND, __A22_NET_90, CCH34, __A22_NET_106, __A22_1__DATA_n, __A22_1__WDORDR, __A22_NET_93, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22027(__A22_1__HIGH0_n, __A22_NET_90, __A22_1__WRD1BP, __A22_1__WRD1B1, __A22_1__WRD2B2, __A22_NET_86, GND, __A22_NET_87, __A22_1__WRD2B3, __A22_NET_88, __A22_NET_89, __A22_NET_89, __A22_1__LOW1_n, p4VDC, SIM_RST, SIM_CLK);
    U74LVC07 U22028(__A22_NET_86, __A22_1__DATA_n, __A22_NET_87, __A22_1__DATA_n, __A22_NET_230, __A22_1__DATA_n, GND, __A22_1__DATA_n, __A22_NET_275, __A22_1__DATA_n, __A22_NET_264, __A22_1__DATA_n, __A22_NET_188, p4VDC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8,10,12
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U22029(__A22_1__DKDAT_n, __A22_NET_93, __A22_1__ORDRBT, __A22_NET_246, WCH34_n, PC15_n, GND, __A22_NET_246, __A22_NET_244, __A22_NET_245, __A22_NET_245, CCH34, __A22_NET_244, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22130(__A22_1__BSYNC_n, __A22_1__RDOUT_n,  ,  ,  ,  , GND,  ,  ,  ,  , __A22_1__DKDATA, __A22_1__DKDAT_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U22131(DKBSNC, __A22_1__BSYNC_n,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U22032(__A22_NET_243, WCH34_n, CHWL01_n, __A22_NET_241, __A22_NET_243, __A22_NET_242, GND, __A22_NET_241, CCH34, __A22_NET_242, WCH34_n, CHWL02_n, __A22_NET_253, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22033(__A22_1__HIGH1_n, __A22_NET_241, __A22_1__HIGH1_n, __A22_NET_254, __A22_1__LOW5_n, __A22_NET_231, GND, __A22_NET_232, __A22_1__HIGH0_n, __A22_NET_248, __A22_1__LOW2_n, __A22_1__WRD1B1, __A22_1__LOW6_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1, 1'b0) U22034(__A22_NET_254, __A22_NET_253, __A22_NET_252, __A22_NET_252, __A22_NET_254, CCH34, GND, WCH34_n, CHWL13_n, __A22_NET_247, __A22_NET_247, __A22_NET_249, __A22_NET_248, p4VDC, SIM_RST, SIM_CLK);
    U74HC4002 U22035(__A22_NET_230, __A22_NET_231, __A22_NET_232, __A22_NET_226, __A22_NET_240,  , GND,  , __A22_NET_276, __A22_NET_236, __A22_NET_271, __A22_NET_274, __A22_NET_275, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U22036(__A22_NET_249, __A22_NET_248, CCH34, __A22_NET_228, WCH34_n, CHWL12_n, GND, __A22_NET_228, __A22_NET_229, __A22_NET_227, __A22_NET_227, CCH34, __A22_NET_229, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22037(__A22_1__HIGH0_n, __A22_NET_227, __A22_1__HIGH0_n, __A22_NET_223, __A22_1__LOW4_n, __A22_NET_240, GND, __A22_NET_276, __A22_1__HIGH0_n, __A22_NET_237, __A22_1__LOW5_n, __A22_NET_226, __A22_1__LOW3_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U22038(__A22_NET_224, WCH34_n, CHWL11_n, __A22_NET_223, __A22_NET_224, __A22_NET_225, GND, __A22_NET_223, CCH34, __A22_NET_225, WCH34_n, CHWL10_n, __A22_NET_238, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1, 1'b0) U22039(__A22_NET_237, __A22_NET_238, __A22_NET_239, __A22_NET_239, __A22_NET_237, CCH34, GND, WCH34_n, CHWL09_n, __A22_NET_233, __A22_NET_233, __A22_NET_235, __A22_NET_234, __A22_NET_54, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U22040(__A22_NET_235, __A22_NET_234, CCH34, __A22_NET_277, WCH34_n, CHWL08_n, GND, __A22_NET_277, __A22_NET_281, __A22_NET_280, __A22_NET_280, CCH34, __A22_NET_281, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22041(__A22_1__HIGH0_n, __A22_NET_234, __A22_1__HIGH0_n, __A22_NET_280, __A22_1__LOW7_n, __A22_NET_271, GND, __A22_NET_274, __A22_1__HIGH1_n, __A22_NET_285, __A22_1__LOW0_n, __A22_NET_236, __A22_1__LOW6_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U22042(__A22_NET_272, WCH34_n, CHWL07_n, __A22_NET_285, __A22_NET_272, __A22_NET_273, GND, __A22_NET_285, CCH34, __A22_NET_273, WCH34_n, CHWL06_n, __A22_NET_288, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1, 1'b0) U22043(__A22_NET_286, __A22_NET_288, __A22_NET_287, __A22_NET_287, __A22_NET_286, CCH34, GND, WCH34_n, CHWL05_n, __A22_NET_282, __A22_NET_282, __A22_NET_283, __A22_NET_284, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22044(__A22_1__HIGH1_n, __A22_NET_286, __A22_1__HIGH1_n, __A22_NET_284, __A22_1__LOW2_n, __A22_NET_266, GND, __A22_NET_260, __A22_1__HIGH1_n, __A22_NET_255, __A22_1__LOW3_n, __A22_NET_263, __A22_1__LOW1_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U22045(__A22_NET_283, __A22_NET_284, CCH34, __A22_NET_267, WCH34_n, CHWL04_n, GND, __A22_NET_267, __A22_NET_256, __A22_NET_255, __A22_NET_255, CCH34, __A22_NET_256, p4VDC, SIM_RST, SIM_CLK);
    U74HC4002 U22046(__A22_NET_264, __A22_NET_263, __A22_NET_266, __A22_NET_260, __A22_NET_262,  , GND,  , __A22_NET_178, __A22_NET_184, __A22_NET_161, __A22_NET_157, __A22_NET_188, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U22047(__A22_NET_257, WCH34_n, CHWL03_n, __A22_NET_258, __A22_NET_257, __A22_NET_259, GND, __A22_NET_258, CCH34, __A22_NET_259, WCH35_n, CHWL16_n, __A22_NET_268, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22048(__A22_1__HIGH1_n, __A22_NET_258, __A22_1__HIGH2_n, __A22_NET_270, __A22_1__LOW0_n, __A22_NET_178, GND, __A22_NET_184, __A22_1__HIGH2_n, __A22_NET_181, __A22_1__LOW1_n, __A22_NET_262, __A22_1__LOW4_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1, 1'b0) U22049(__A22_NET_270, __A22_NET_268, __A22_NET_269, __A22_NET_269, __A22_NET_270, CCH35, GND, WCH35_n, CHWL14_n, __A22_NET_183, __A22_NET_183, __A22_NET_182, __A22_NET_181, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U22050(__A22_NET_182, __A22_NET_181, CCH35, __A22_NET_177, WCH35_n, CHWL13_n, GND, __A22_NET_177, __A22_NET_176, __A22_NET_175, __A22_NET_175, CCH35, __A22_NET_176, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22051(__A22_1__HIGH2_n, __A22_NET_175, __A22_1__HIGH2_n, __A22_NET_191, __A22_1__LOW3_n, __A22_NET_157, GND, __A22_NET_165, __A22_1__HIGH2_n, __A22_NET_185, __A22_1__LOW4_n, __A22_NET_161, __A22_1__LOW2_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U22052(__A22_NET_189, WCH35_n, CHWL12_n, __A22_NET_191, __A22_NET_189, __A22_NET_190, GND, __A22_NET_191, CCH35, __A22_NET_190, WCH35_n, CHWL11_n, __A22_NET_186, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1, 1'b0) U22053(__A22_NET_185, __A22_NET_186, __A22_NET_187, __A22_NET_187, __A22_NET_185, CCH35, GND, WCH35_n, CHWL10_n, __A22_NET_158, __A22_NET_158, __A22_NET_160, __A22_NET_159, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U22054(__A22_NET_160, __A22_NET_159, CCH35, __A22_NET_155, WCH35_n, CHWL09_n, GND, __A22_NET_155, __A22_NET_156, __A22_NET_154, __A22_NET_154, CCH35, __A22_NET_156, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22055(__A22_1__HIGH2_n, __A22_NET_159, __A22_1__HIGH2_n, __A22_NET_154, __A22_1__LOW6_n, __A22_NET_169, GND, __A22_NET_168, __A22_1__HIGH2_n, __A22_NET_174, __A22_1__LOW7_n, __A22_NET_162, __A22_1__LOW5_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC4002 U22056(__A22_NET_164, __A22_NET_165, __A22_NET_162, __A22_NET_169, __A22_NET_168,  , GND,  , __A22_NET_216, __A22_NET_215, __A22_NET_196, __A22_NET_195, __A22_NET_214, p4VDC, SIM_RST, SIM_CLK);
    U74LVC07 U22057(__A22_NET_164, __A22_1__DATA_n, __A22_NET_214, __A22_1__DATA_n, __A22_NET_203, __A22_1__DATA_n, GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U22058(__A22_NET_173, WCH35_n, CHWL08_n, __A22_NET_174, __A22_NET_173, __A22_NET_172, GND, __A22_NET_174, CCH35, __A22_NET_172, WCH35_n, CHWL07_n, __A22_NET_163, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1, 1'b0) U22059(__A22_NET_171, __A22_NET_163, __A22_NET_170, __A22_NET_170, __A22_NET_171, CCH35, GND, WCH35_n, CHWL06_n, __A22_NET_210, __A22_NET_210, __A22_NET_211, __A22_NET_212, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22060(__A22_1__HIGH3_n, __A22_NET_171, __A22_1__HIGH3_n, __A22_NET_212, __A22_1__LOW1_n, __A22_NET_215, GND, __A22_NET_196, __A22_1__HIGH3_n, __A22_NET_209, __A22_1__LOW2_n, __A22_NET_216, __A22_1__LOW0_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U22061(__A22_NET_211, __A22_NET_212, CCH35, __A22_NET_208, WCH35_n, CHWL05_n, GND, __A22_NET_208, __A22_NET_207, __A22_NET_209, __A22_NET_209, CCH35, __A22_NET_207, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U22062(__A22_NET_220, WCH35_n, CHWL04_n, __A22_NET_222, __A22_NET_220, __A22_NET_221, GND, __A22_NET_222, CCH35, __A22_NET_221, WCH35_n, CHWL03_n, __A22_NET_218, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22063(__A22_1__HIGH3_n, __A22_NET_222, __A22_1__HIGH3_n, __A22_NET_197, __A22_1__LOW4_n, __A22_1__WRD2B3, GND, __A22_1__WRD2B2, __A22_1__HIGH3_n, __A22_NET_192, __A22_1__LOW5_n, __A22_NET_195, __A22_1__LOW3_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1, 1'b0) U22064(__A22_NET_197, __A22_NET_218, __A22_NET_219, __A22_NET_219, __A22_NET_197, CCH35, GND, WCH35_n, CHWL02_n, __A22_NET_199, __A22_NET_199, __A22_NET_198, __A22_NET_192, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U22065(__A22_NET_198, __A22_NET_192, CCH35, __A22_NET_193, WCH35_n, CHWL01_n, GND, __A22_NET_193, __A22_NET_205, __A22_NET_204, __A22_NET_204, CCH35, __A22_NET_205, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22066(__A22_1__HIGH3_n, __A22_NET_204, __A22_1__HIGH3_n, __A22_NET_200, __A22_1__LOW7_n, __A22_NET_202, GND,  ,  ,  ,  , __A22_NET_194, __A22_1__LOW6_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U22067(__A22_NET_206, WCH35_n, PC15_n, __A22_NET_200, __A22_NET_206, __A22_NET_201, GND, __A22_NET_200, CCH35, __A22_NET_201, __A22_NET_194, __A22_NET_202, __A22_NET_203, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22068(__A22_1__BSYNC_n, __A22_1__RDOUT_n, __A22_1__HIGH1_n, __A22_NET_245, __A22_1__LOW7_n, __A22_1__WRD1BP, GND,  ,  ,  ,  , __A22_1__DKDATB, __A22_1__DKDAT_n, p4VDC, SIM_RST, SIM_CLK);
endmodule