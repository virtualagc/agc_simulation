`timescale 1ns/1ps

module crosspoint_nqi(VCC, GND, SIM_RST, GOJAM, T01, T01_n, T02_n, T03_n, T04_n, T05_n, T06_n, T07_n, T08_n, T09_n, T10_n, T11_n, T12, T12_n, T12USE_n, STD2, BR1, BR1_n, BR2, BR2_n, BR12B_n, BR1B2_n, BRDIF_n, S11, S12, INCSET_n, INKL_n, MONPCH, MONWBK, ADS0, CCS0, CCS0_n, CHINC_n, DAS0, DAS0_n, DAS1, DAS1_n, DV1, DV1_n, DV4, DV4_n, DIV_n, DXCH0, FETCH0, FETCH0_n, GOJ1, GOJ1_n, INOUT, INOUT_n, MASK0, MASK0_n, MP0, MP3, MP3_n, MSU0, MSU0_n, NDX0_n, PRINC, QXCH0_n, RAND0, READ0, ROR0, RSM3, RSM3_n, RUPT0, RXOR0, RXOR0_n, SHANC_n, SHIFT, SHIFT_n, STFET1_n, TC0, TC0_n, TCF0, TCSAJ3_n, TS0, TS0_n, WAND0, WOR0, IC1, IC2, IC2_n, IC3, IC4, IC5, IC5_n, IC8_n, IC9, IC10, IC10_n, IC11_n, IC12, IC12_n, IC13, IC14, IC15_n, IC16, IC16_n, C24A, C25A, C26A, C27A, C30A, C37P, C40P, C41P, C42P, C43P, C44P, XT0_n, XT2_n, XT3_n, XT4_n, XT5_n, XT6_n, YB0_n, YT0_n, n4XP5, n5XP9, n5XP11, n10XP6, A2X_n, CI_n, PINC, DVST, MONEX_n, NDR100_n, NISQ, PTWOX, R6, RA_n, RAD, RB_n, RC_n, RG_n, RL_n, RL10BB, RQ_n, RSTSTG, RU_n, RZ_n, SCAD, SCAD_n, ST2_n, TMZ_n, TOV_n, TPZG_n, TSGN_n, TSUDO_n, U2BBK, WA_n, WB_n, WG_n, WL_n, WS_n, WY_n, WY12_n, WYD_n, WZ_n, DV4B1B, TRSM, OCTAD2, n2XP7, n2XP8, n3XP6, n5XP12, n5XP15, n5XP21, n6XP8, n7XP4, n7XP9, n9XP5, n10XP1, n10XP8, n11XP2);
    input wire SIM_RST;
    inout wire A2X_n;
    input wire ADS0;
    input wire BR1;
    input wire BR12B_n;
    input wire BR1B2_n;
    input wire BR1_n;
    input wire BR2;
    input wire BR2_n;
    input wire BRDIF_n;
    input wire C24A;
    input wire C25A;
    input wire C26A;
    input wire C27A;
    input wire C30A;
    input wire C37P;
    input wire C40P;
    input wire C41P;
    input wire C42P;
    input wire C43P;
    input wire C44P;
    input wire CCS0;
    input wire CCS0_n;
    input wire CHINC_n;
    inout wire CI_n;
    input wire DAS0;
    input wire DAS0_n;
    input wire DAS1;
    input wire DAS1_n;
    input wire DIV_n;
    input wire DV1;
    input wire DV1_n;
    input wire DV4;
    output wire DV4B1B;
    input wire DV4_n;
    output wire DVST;
    input wire DXCH0;
    input wire FETCH0;
    input wire FETCH0_n;
    input wire GND;
    input wire GOJ1;
    input wire GOJ1_n;
    input wire GOJAM;
    input wire IC1;
    input wire IC10;
    input wire IC10_n;
    input wire IC11_n;
    input wire IC12;
    input wire IC12_n;
    input wire IC13;
    input wire IC14;
    input wire IC15_n;
    input wire IC16;
    input wire IC16_n;
    input wire IC2;
    input wire IC2_n;
    input wire IC3;
    input wire IC4;
    input wire IC5;
    input wire IC5_n;
    input wire IC8_n;
    input wire IC9;
    input wire INCSET_n;
    input wire INKL_n;
    input wire INOUT;
    input wire INOUT_n;
    input wire MASK0;
    input wire MASK0_n;
    inout wire MONEX_n;
    input wire MONPCH;
    input wire MONWBK;
    input wire MP0;
    input wire MP3;
    input wire MP3_n;
    input wire MSU0;
    input wire MSU0_n;
    output wire NDR100_n;
    input wire NDX0_n;
    wire NET_195;
    wire NET_196;
    wire NET_197;
    wire NET_198;
    wire NET_199;
    wire NET_200;
    wire NET_201;
    wire NET_202;
    wire NET_203;
    wire NET_204;
    wire NET_205;
    wire NET_208;
    wire NET_209;
    wire NET_211;
    wire NET_212;
    wire NET_213;
    wire NET_214;
    wire NET_216;
    wire NET_217;
    wire NET_218;
    wire NET_219;
    wire NET_220;
    wire NET_221;
    wire NET_222;
    wire NET_225;
    wire NET_226;
    wire NET_227;
    wire NET_228;
    wire NET_229;
    wire NET_230;
    wire NET_231;
    wire NET_232;
    wire NET_233;
    wire NET_234;
    wire NET_235;
    wire NET_236;
    wire NET_237;
    wire NET_238;
    wire NET_239;
    wire NET_240;
    wire NET_241;
    wire NET_242;
    wire NET_243;
    wire NET_244;
    wire NET_245;
    wire NET_246;
    wire NET_247;
    wire NET_248;
    wire NET_249;
    wire NET_250;
    wire NET_251;
    wire NET_252;
    wire NET_253;
    wire NET_254;
    wire NET_255;
    wire NET_256;
    wire NET_258;
    wire NET_259;
    wire NET_260;
    wire NET_261;
    wire NET_262;
    wire NET_263;
    wire NET_264;
    wire NET_265;
    wire NET_266;
    wire NET_267;
    wire NET_268;
    wire NET_269;
    wire NET_270;
    wire NET_271;
    wire NET_272;
    wire NET_273;
    wire NET_274;
    wire NET_275;
    wire NET_276;
    wire NET_277;
    wire NET_278;
    wire NET_279;
    wire NET_280;
    wire NET_281;
    wire NET_282;
    wire NET_283;
    wire NET_284;
    wire NET_285;
    wire NET_286;
    wire NET_287;
    wire NET_288;
    wire NET_289;
    wire NET_290;
    wire NET_291;
    wire NET_292;
    wire NET_294;
    wire NET_295;
    wire NET_296;
    wire NET_297;
    wire NET_298;
    wire NET_299;
    wire NET_300;
    wire NET_302;
    wire NET_303;
    wire NET_304;
    wire NET_305;
    wire NET_306;
    wire NET_308;
    wire NET_309;
    wire NET_310;
    wire NET_311;
    wire NET_312;
    wire NET_313;
    wire NET_314;
    wire NET_315;
    wire NET_316;
    wire NET_317;
    wire NET_318;
    wire NET_320;
    wire NET_321;
    wire NET_322;
    wire NET_323;
    wire NET_324;
    wire NET_325;
    wire NET_327;
    wire NET_328;
    wire NET_329;
    wire NET_330;
    wire NET_331;
    wire NET_332;
    wire NET_333;
    wire NET_334;
    wire NET_335;
    wire NET_337;
    wire NET_339;
    wire NET_341;
    wire NET_342;
    wire NET_343;
    wire NET_344;
    wire NET_345;
    wire NET_346;
    wire NET_347;
    wire NET_348;
    wire NET_349;
    wire NET_350;
    wire NET_351;
    wire NET_352;
    wire NET_353;
    wire NET_354;
    wire NET_355;
    wire NET_356;
    wire NET_357;
    wire NET_358;
    wire NET_359;
    wire NET_360;
    wire NET_361;
    wire NET_362;
    wire NET_363;
    wire NET_364;
    wire NET_365;
    wire NET_366;
    wire NET_367;
    wire NET_368;
    wire NET_369;
    wire NET_370;
    wire NET_371;
    wire NET_372;
    wire NET_373;
    output wire NISQ;
    output wire OCTAD2;
    output wire PINC;
    input wire PRINC;
    output wire PTWOX;
    input wire QXCH0_n;
    output wire R6;
    output wire RAD;
    input wire RAND0;
    inout wire RA_n;
    inout wire RB_n;
    inout wire RC_n;
    input wire READ0;
    inout wire RG_n;
    output wire RL10BB;
    inout wire RL_n;
    input wire ROR0;
    output wire RQ_n;
    input wire RSM3;
    input wire RSM3_n;
    output wire RSTSTG;
    input wire RUPT0;
    inout wire RU_n;
    input wire RXOR0;
    input wire RXOR0_n;
    inout wire RZ_n;
    input wire S11;
    input wire S12;
    inout wire SCAD;
    output wire SCAD_n;
    input wire SHANC_n;
    input wire SHIFT;
    input wire SHIFT_n;
    inout wire ST2_n;
    input wire STD2;
    input wire STFET1_n;
    input wire T01;
    input wire T01_n;
    input wire T02_n;
    input wire T03_n;
    input wire T04_n;
    input wire T05_n;
    input wire T06_n;
    input wire T07_n;
    input wire T08_n;
    input wire T09_n;
    input wire T10_n;
    input wire T11_n;
    input wire T12;
    input wire T12USE_n;
    input wire T12_n;
    input wire TC0;
    input wire TC0_n;
    input wire TCF0;
    input wire TCSAJ3_n;
    inout wire TMZ_n;
    inout wire TOV_n;
    output wire TPZG_n;
    output wire TRSM;
    input wire TS0;
    input wire TS0_n;
    output wire TSGN_n;
    output wire TSUDO_n;
    output wire U2BBK;
    input wire VCC;
    input wire WAND0;
    inout wire WA_n;
    inout wire WB_n;
    inout wire WG_n;
    inout wire WL_n;
    input wire WOR0;
    inout wire WS_n;
    inout wire WY12_n;
    inout wire WYD_n;
    inout wire WY_n;
    inout wire WZ_n;
    input wire XT0_n;
    input wire XT2_n;
    input wire XT3_n;
    input wire XT4_n;
    input wire XT5_n;
    input wire XT6_n;
    input wire YB0_n;
    input wire YT0_n;
    wire __A05_1__10XP7;
    wire __A05_1__3XP5;
    wire __A05_1__8XP12;
    wire __A05_1__8XP15;
    wire __A05_1__8XP3;
    wire __A05_1__DV1B1B;
    wire __A05_1__GHNHC;
    wire __A05_1__MNISQ;
    wire __A05_1__NISQ_n;
    wire __A05_1__PARTC;
    wire __A05_1__PINC_n;
    wire __A05_1__RSTRT;
    wire __A05_2__10XP10;
    wire __A05_2__11XP6;
    wire __A05_2__5XP13;
    wire __A05_2__5XP19;
    wire __A05_2__6XP2;
    wire __A05_2__6XP7;
    wire __A05_2__OCTAD3;
    wire __A05_2__OCTAD4;
    wire __A05_2__OCTAD5;
    wire __A05_2__OCTAD6;
    wire __A05_2__RSCT;
    wire __A05_2__Z15_n;
    wire __A05_2__Z16_n;
    output wire n10XP1;
    output wire n10XP6;
    output wire n10XP8;
    output wire n11XP2;
    output wire n2XP7;
    output wire n2XP8;
    output wire n3XP6;
    input wire n4XP5;
    input wire n5XP11;
    output wire n5XP12;
    output wire n5XP15;
    output wire n5XP21;
    output wire n5XP9;
    output wire n6XP8;
    output wire n7XP4;
    output wire n7XP9;
    output wire n9XP5;

    pullup R5001(NET_216);
    pullup R5002(NET_311);
    pullup R5003(NET_313);
    pullup R5004(RL_n);
    pullup R5005(RA_n);
    pullup R5006(WY_n);
    pullup R5007(WY12_n);
    pullup R5008(SCAD);
    pullup R5009(NET_329);
    pullup R5010(NET_331);
    pullup R5011(TMZ_n);
    U74HC27 U5001(IC10, IC3, TC0, TCF0, IC4, NET_248, GND, NET_247, IC2, IC3, RSM3, NET_250, IC2, VCC, SIM_RST);
    U74HC02 U5002(NET_249, STD2, IC2, NET_271, T01_n, NET_250, GND, T01_n, NET_249, NET_252, IC10_n, T01_n, NET_253, VCC, SIM_RST);
    U74HC02 U5003(NET_268, T01_n, NET_248, NET_251, T02_n, NET_247, GND, T08_n, CCS0_n, NET_212, T02_n, MP3_n, n2XP7, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U5004(T02_n, STD2, n10XP6, __A05_1__10XP7, NET_253, NET_256, GND, NET_260, NET_252, n3XP6, NET_243, DVST, DIV_n, VCC, SIM_RST);
    U74LVC07 U5005(NET_256, MONEX_n, NET_260, RZ_n, NET_261, RB_n, GND, RA_n, NET_258, WA_n, NET_246, RL_n, NET_240, VCC, SIM_RST);
    U74HC27 U5006(NET_251, __A05_1__8XP15, NET_241, NET_244, __A05_1__8XP12, NET_240, GND, __A05_1__PARTC, INKL_n, SHIFT, MONPCH, __A05_1__NISQ_n, n2XP7, VCC, SIM_RST);
    U74HC02 U5007(__A05_1__3XP5, T03_n, IC2_n, NET_276, T01_n, IC15_n, GND, NET_276, NET_259, NET_258, T03_n, TC0_n, n3XP6, VCC, SIM_RST);
    U74HC02 U5008(NET_259, T04_n, IC2_n, NET_245, T02_n, IC15_n, GND, NET_245, NET_275, TPZG_n, T04_n, DAS0_n, NET_241, VCC, SIM_RST);
    U74HC02 #(1, 0, 0, 0) U5009(NET_246, NET_241, NET_242, NET_242, T04_n, MASK0_n, GND, MP3_n, T10_n, NET_244, T05_n, IC2_n, NET_243, VCC, SIM_RST);
    U74HC02 U5010(NET_275, T05_n, NET_255, NET_254, NET_276, NET_275, GND, T05_n, DAS0_n, n5XP12, T06_n, RSM3_n, NET_280, VCC, SIM_RST);
    U74HC27 U5011(__A05_1__PARTC, PRINC, NET_275, NET_276, n7XP9, TSGN_n, GND, NET_281, n9XP5, NET_276, NET_280, NET_255, CCS0, VCC, SIM_RST);
    U74LVC07 U5012(NET_254, TMZ_n, NET_281, WG_n, NET_278, RG_n, GND, RC_n, NET_279, A2X_n, NET_263, WY_n, NET_265, VCC, SIM_RST);
    U74HC02 U5013(NET_264, T06_n, DAS0_n, NET_277, T06_n, MSU0_n, GND, NET_242, NET_277, NET_279, T07_n, DAS0_n, NET_267, VCC, SIM_RST);
    U74HC27 #(0, 1, 1) U5014(NET_275, NET_262, NET_262, NET_264, NET_277, NET_263, GND, NET_265, NET_262, NET_277, NET_264, NET_278, NET_264, VCC, SIM_RST);
    U74HC4002 U5015(NET_261, NET_268, __A05_1__3XP5, NET_267, NET_280, NET_266, GND, NET_269, IC3, RSM3, MP3, IC16, TSUDO_n, VCC, SIM_RST);
    U74HC02 U5016(n7XP9, T07_n, MSU0_n, NET_262, T07_n, IC2_n, GND, T07_n, CCS0_n, NET_274, NET_203, NET_195, NET_204, VCC, SIM_RST);
    U74HC27 #(0, 0, 1) U5017(NET_277, NET_271, __A05_1__8XP3, NET_274, n4XP5, NET_272, GND, NET_270, n4XP5, NET_274, NET_271, NET_273, n10XP6, VCC, SIM_RST);
    U74LVC07 U5018(NET_273, CI_n, NET_272, RZ_n, NET_270, WY12_n, GND, WZ_n, NET_205, RB_n, NET_204, WB_n, NET_213, VCC, SIM_RST);
    U74HC27 #(0, 0, 1) U5019(CCS0_n, T07_n, BR1_n, CCS0_n, T07_n, PTWOX, GND, NET_205, __A05_1__3XP5, NET_197, NET_212, n7XP4, BR2_n, VCC, SIM_RST);
    U74HC27 U5020(INKL_n, FETCH0, NET_212, NET_209, n9XP5, NET_199, GND, NET_211, IC2, IC4, DXCH0, NET_203, T08_n, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U5021(RAD, TSUDO_n, T08_n, NET_213, RAD, NET_200, GND, T08_n, NET_214, __A05_1__8XP15, T08_n, NET_208, __A05_1__8XP3, VCC, SIM_RST);
    U74HC04 U5022(IC16, NET_214, NET_289, RQ_n, MP3, NET_299, GND, SCAD_n, SCAD, NDR100_n, NET_292, NET_335, NET_328, VCC, SIM_RST);
    U74HC02 U5023(NET_208, MP0, IC1, NET_209, T08_n, NET_211, GND, T08_n, NET_198, NET_200, T08_n, GOJ1_n, __A05_1__RSTRT, VCC, SIM_RST);
    U74LVC07 U5024(NET_199, RU_n, NET_202, RA_n, NET_201, ST2_n, GND, WY_n, NET_233, RC_n, NET_237, WA_n, NET_221, VCC, SIM_RST);
    U74HC27 U5025(DXCH0, GOJ1, T08_n, BR2, T10_n, n10XP6, GND, NET_235, IC1, IC10, RUPT0, NET_198, DAS0, VCC, SIM_RST);
    U74HC02 U5026(__A05_1__8XP12, T08_n, DAS0_n, NET_197, T08_n, TCSAJ3_n, GND, T09_n, NET_196, NET_195, IC2, __A05_1__DV1B1B, NET_196, VCC, SIM_RST);
    U74HC02 U5027(n9XP5, T09_n, DAS0_n, NET_231, T09_n, MASK0_n, GND, NET_231, NET_232, NET_202, T10_n, T08_n, NET_229, VCC, SIM_RST);
    U74HC02 U5028(NET_201, NET_197, NET_229, n10XP1, NET_235, T10_n, GND, T10_n, NET_230, NET_232, DAS0, NET_239, NET_230, VCC, SIM_RST);
    U74HC27 #(1, 0, 1) U5029(NET_229, NET_231, T10_n, DAS0_n, BR1B2_n, n10XP8, GND, NET_221, NET_195, NET_220, n5XP11, NET_233, NET_232, VCC, SIM_RST);
    U74HC02 U5030(NET_239, MSU0_n, BR1_n, __A05_1__10XP7, T10_n, NET_234, GND, NET_239, NET_238, NET_234, BR12B_n, DAS0_n, NET_238, VCC, SIM_RST);
    U74HC02 U5031(n11XP2, T11_n, MSU0_n, NET_236, T10_n, MASK0_n, GND, NET_231, NET_236, NET_237, T10_n, NET_222, NET_220, VCC, SIM_RST);
    U74HC02 U5032(NET_222, MSU0, IC14, NET_227, INCSET_n, NET_216, GND, GOJAM, __A05_1__GHNHC, NET_228, NET_228, T01, __A05_1__GHNHC, VCC, SIM_RST);
    U74HC4002 U5033(NET_218, C24A, C25A, C26A, C27A, NET_226, GND, NET_225, C30A, C37P, C40P, C41P, NET_217, VCC, SIM_RST);
    U74HC27 #(0, 0, 1) U5034(C42P, C43P, IC12, DAS0, DAS1, NET_354, GND, NET_350, RL10BB, NET_310, __A05_2__RSCT, NET_219, C44P, VCC, SIM_RST);
    U74LVC07 U5035(NET_218, NET_216, NET_217, NET_216, NET_219, NET_216, GND, NET_311, NET_354, NET_311, NET_353, WS_n, NET_350, VCC, SIM_RST);
    U74HC02 U5036(__A05_1__PINC_n, NET_227, PINC, PINC, __A05_1__PINC_n, T12, GND, T01_n, NET_311, RL10BB, T01_n, FETCH0_n, R6, VCC, SIM_RST);
    U74HC4002 U5037(NET_353, IC9, DXCH0, PRINC, INOUT, NET_352, GND, NET_351, YB0_n, YT0_n, S12, S11, NET_292, VCC, SIM_RST);
    U74HC02 U5038(NET_310, T01_n, CHINC_n, NET_286, T03_n, NET_313, GND, IC5, MP0, NET_355, T03_n, IC8_n, NET_312, VCC, SIM_RST);
    U74HC27 #(0, 0, 1) U5039(T01_n, MONPCH, TS0, DAS0, MASK0, NET_358, GND, NET_356, NET_286, NET_312, NET_289, __A05_2__RSCT, INKL_n, VCC, SIM_RST);
    wire U5040_3_NC;
    wire U5040_4_NC;
    wire U5040_5_NC;
    wire U5040_6_NC;
    wire U5040_8_NC;
    wire U5040_9_NC;
    wire U5040_10_NC;
    wire U5040_11_NC;
    U74HC27 #(1, 0, 0) U5040(NET_287, NET_290, U5040_3_NC, U5040_4_NC, U5040_5_NC, U5040_6_NC, GND, U5040_8_NC, U5040_9_NC, U5040_10_NC, U5040_11_NC, NET_357, __A05_2__6XP2, VCC, SIM_RST);
    U74LVC07 U5041(NET_356, WB_n, NET_357, WB_n, NET_358, NET_313, GND, NET_313, NET_355, RL_n, NET_345, RA_n, NET_346, VCC, SIM_RST);
    U74HC02 U5042(n2XP8, T02_n, FETCH0_n, NET_289, T03_n, QXCH0_n, GND, T04_n, DV1_n, NET_288, T04_n, NET_291, NET_287, VCC, SIM_RST);
    U74HC27 U5043(NET_312, NET_288, DV1, INOUT, IC2, NET_291, GND, NET_344, NET_290, NET_285, n5XP9, NET_345, __A05_2__11XP6, VCC, SIM_RST);
    U74HC02 U5044(NET_346, NET_286, __A05_2__6XP2, TRSM, T05_n, NDX0_n, GND, IC12_n, T05_n, NET_290, DAS1_n, T05_n, NET_285, VCC, SIM_RST);
    U74HC27 #(0, 0, 1) U5045(__A05_2__5XP13, n5XP15, DAS1, PRINC, __A05_1__PARTC, NET_282, GND, NET_349, NET_283, n2XP8, __A05_2__10XP10, NET_343, NET_297, VCC, SIM_RST);
    U74LVC07 U5046(NET_344, RG_n, NET_343, RG_n, NET_349, WY_n, GND, A2X_n, NET_347, CI_n, NET_348, WY12_n, NET_371, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U5047(NET_283, NET_282, T05_n, NET_347, NET_285, __A05_2__10XP10, GND, SHIFT_n, T05_n, n5XP9, SHANC_n, T05_n, NET_284, VCC, SIM_RST);
    U74HC27 U5048(NET_284, NET_298, YT0_n, YB0_n, XT0_n, NET_372, GND, NET_296, RAND0, WAND0, NET_328, NET_348, NET_300, VCC, SIM_RST);
    U74HC02 U5049(__A05_2__5XP13, IC8_n, T05_n, n5XP15, QXCH0_n, T05_n, GND, CHINC_n, T05_n, n5XP21, IC5_n, T05_n, NET_297, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U5050(NET_298, IC16_n, T05_n, NET_300, NET_299, T05_n, GND, NET_298, NET_300, NET_371, S11, S12, NET_373, VCC, SIM_RST);
    U74LVC07 U5051(NET_370, RB_n, NET_369, RZ_n, NET_373, SCAD, GND, SCAD, NET_372, RC_n, NET_362, NET_329, NET_360, VCC, SIM_RST);
    U74HC02 U5052(NET_370, __A05_2__5XP19, NET_298, NET_369, __A05_2__6XP7, NET_300, GND, XT2_n, NDR100_n, OCTAD2, NDR100_n, XT3_n, __A05_2__OCTAD3, VCC, SIM_RST);
    U74HC02 U5053(__A05_2__OCTAD4, NDR100_n, XT4_n, __A05_2__OCTAD5, NDR100_n, XT5_n, GND, NDR100_n, XT6_n, __A05_2__OCTAD6, BR1_n, DV1_n, NET_328, VCC, SIM_RST);
    U74HC02 U5054(NET_295, NET_296, T05_n, __A05_2__5XP19, T05_n, NET_294, GND, DV1_n, BR1, __A05_1__DV1B1B, TS0_n, BRDIF_n, NET_330, VCC, SIM_RST);
    U74HC4002 #(0, 1) U5055(NET_362, NET_295, NET_332, NET_324, NET_323, NET_361, GND, NET_363, __A05_2__5XP13, NET_308, NET_339, NET_317, NET_337, VCC, SIM_RST);
    U74HC27 U5056(ROR0, __A05_1__DV1B1B, IC2, IC5, READ0, NET_360, GND, NET_364, IC2, IC3, TS0, NET_294, WOR0, VCC, SIM_RST);
    U74HC02 #(0, 0, 0, 1) U5057(NET_359, NET_330, DV4, NET_333, NET_329, T05_n, GND, NET_335, T05_n, NET_334, NET_333, NET_332, NET_367, VCC, SIM_RST);
    U74LVC07 U5058(NET_359, NET_329, NET_368, __A05_2__Z16_n, NET_367, WA_n, GND, NET_331, NET_364, NET_331, NET_365, WZ_n, NET_366, VCC, SIM_RST);
    U74HC04 #(0, 1, 0, 0, 0, 0) U5059(NET_334, NET_368, NET_327, NET_366, NET_332, NET_342, GND, NET_322, NET_324, NISQ, __A05_1__NISQ_n, __A05_1__MNISQ, __A05_1__NISQ_n, VCC, SIM_RST);
    U74HC02 U5060(NET_365, IC16, MP3, NET_327, T06_n, NET_331, GND, T06_n, DAS1_n, n6XP8, n6XP8, __A05_2__6XP7, NET_306, VCC, SIM_RST);
    U74LVC07 U5061(NET_306, TOV_n, NET_303, RU_n, NET_302, RU_n, GND, WB_n, NET_304, RG_n, NET_314, TSGN_n, NET_341, VCC, SIM_RST);
    U74HC02 U5062(__A05_2__6XP7, DV4_n, T06_n, NET_316, T07_n, NET_305, GND, T07_n, STFET1_n, NET_315, T08_n, DV4_n, RSTSTG, VCC, SIM_RST);
    U74HC27 U5063(NET_327, n6XP8, NET_309, NET_339, NET_308, NET_302, GND, __A05_2__6XP2, T06_n, RXOR0, INOUT_n, NET_303, n5XP11, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U5064(IC13, IC14, NET_316, NET_339, NET_309, NET_304, GND, NET_314, NET_316, NET_315, NET_323, NET_305, DV1, VCC, SIM_RST);
    U74HC27 U5065(T08_n, MONWBK, IC2, IC14, DV1, NET_321, GND, NET_318, DV4B1B, IC4, NET_320, U2BBK, STFET1_n, VCC, SIM_RST);
    U74HC02 U5066(NET_341, RSTSTG, n5XP9, NET_332, T09_n, NET_335, GND, T09_n, DV4_n, NET_339, T09_n, DAS1_n, NET_324, VCC, SIM_RST);
    wire U5067_10_NC;
    wire U5067_11_NC;
    wire U5067_12_NC;
    wire U5067_13_NC;
    U74LVC07 U5067(NET_342, __A05_2__Z15_n, NET_337, WL_n, NET_322, TMZ_n, GND, WYD_n, NET_325, U5067_10_NC, U5067_11_NC, U5067_12_NC, U5067_13_NC, VCC, SIM_RST);
    wire U5068_4_NC;
    wire U5068_5_NC;
    wire U5068_6_NC;
    U74HC02 U5068(NET_309, T10_n, NET_321, U5068_4_NC, U5068_5_NC, U5068_6_NC, GND, T10_n, IC11_n, __A05_2__10XP10, T10_n, NET_318, NET_317, VCC, SIM_RST);
    wire U5069_8_NC;
    wire U5069_9_NC;
    wire U5069_10_NC;
    wire U5069_11_NC;
    U74HC27 U5069(DAS1_n, ADS0, T12_n, T12USE_n, DV1_n, NET_308, GND, U5069_8_NC, U5069_9_NC, U5069_10_NC, U5069_11_NC, NET_320, BR2, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U5070(DV4B1B, DV4_n, BR1, __A05_2__11XP6, T11_n, DV1_n, GND, n5XP9, __A05_2__11XP6, NET_325, T11_n, RXOR0_n, NET_323, VCC, SIM_RST);
endmodule