`timescale 1ns/1ps

module crosspoint_ii(VCC, GND, SIM_RST, GOJAM, T01, T01_n, T02, T02_n, T03, T03_n, T04, T04_n, T05, T06, T06_n, T07, T07_n, T08, T08_n, T09, T10, T10_n, T11, T11_n, T12, T12USE_n, PHS4_n, ST2_n, BR1, BR1_n, BR2_n, BR1B2_n, BR12B_n, BR1B2B, BR1B2B_n, INKL, AD0, ADS0, AUG0_n, CCS0, CCS0_n, CDUSTB_n, DAS0, DAS1, DAS1_n, DCA0, DCS0, DIM0_n, DINC, DINC_n, DV1376, DV1376_n, DV376_n, DV4_n, DV4B1B, DXCH0, FETCH1, INCR0, INOTLD, MASK0, MCDU, MINC, MP0T10, MP1, MP1_n, MP3_n, MSU0, NDXX1_n, PCDU, PINC, PRINC, RAND0, RUPT0, RUPT1, SHIFT, STFET1_n, SU0, WAND0, IC6, IC7, IC9, IC11, IC17, B15X, DIVSTG, PTWOX, R6, R15, RADRG, RADRZ, RBSQ, RRPA, STBE, STBF, TL15, L01_n, L02A_n, L15A_n, MON_n, MONPCH, n8PP4, n1XP10, n2XP3, n2XP5, n2XP7, n2XP8, n3XP2, n3XP6, n3XP7, n4XP11, n5XP4, n5XP12, n5XP15, n5XP21, n5XP28, n6XP5, n6XP8, n7XP4, n7XP9, n7XP19, n8XP6, n9XP1, n9XP5, n10XP1, n10XP8, n11XP2, EXT, MONEX_n, ST1, ST2, TSGU_n, n7XP14);
    input wire SIM_RST;
    input wire AD0;
    input wire ADS0;
    input wire AUG0_n;
    input wire B15X;
    input wire BR1;
    input wire BR12B_n;
    input wire BR1B2B;
    input wire BR1B2B_n;
    input wire BR1B2_n;
    input wire BR1_n;
    input wire BR2_n;
    input wire CCS0;
    input wire CCS0_n;
    input wire CDUSTB_n;
    input wire DAS0;
    input wire DAS1;
    input wire DAS1_n;
    input wire DCA0;
    input wire DCS0;
    input wire DIM0_n;
    input wire DINC;
    input wire DINC_n;
    input wire DIVSTG;
    input wire DV1376;
    input wire DV1376_n;
    input wire DV376_n;
    input wire DV4B1B;
    input wire DV4_n;
    input wire DXCH0;
    output wire EXT;
    input wire FETCH1;
    input wire GND;
    input wire GOJAM;
    input wire IC11;
    input wire IC17;
    input wire IC6;
    input wire IC7;
    input wire IC9;
    input wire INCR0;
    input wire INKL;
    input wire INOTLD;
    input wire L01_n;
    input wire L02A_n;
    input wire L15A_n;
    input wire MASK0;
    input wire MCDU;
    input wire MINC;
    inout wire MONEX_n;
    input wire MONPCH;
    input wire MON_n;
    input wire MP0T10;
    input wire MP1;
    input wire MP1_n;
    input wire MP3_n;
    input wire MSU0;
    input wire NDXX1_n;
    wire NET_181;
    wire NET_182;
    wire NET_183;
    wire NET_184;
    wire NET_185;
    wire NET_187;
    wire NET_188;
    wire NET_189;
    wire NET_190;
    wire NET_191;
    wire NET_193;
    wire NET_194;
    wire NET_195;
    wire NET_196;
    wire NET_199;
    wire NET_200;
    wire NET_201;
    wire NET_202;
    wire NET_203;
    wire NET_204;
    wire NET_205;
    wire NET_206;
    wire NET_207;
    wire NET_208;
    wire NET_209;
    wire NET_210;
    wire NET_212;
    wire NET_213;
    wire NET_214;
    wire NET_215;
    wire NET_216;
    wire NET_217;
    wire NET_218;
    wire NET_219;
    wire NET_220;
    wire NET_222;
    wire NET_223;
    wire NET_224;
    wire NET_227;
    wire NET_229;
    wire NET_230;
    wire NET_231;
    wire NET_232;
    wire NET_233;
    wire NET_235;
    wire NET_236;
    wire NET_238;
    wire NET_239;
    wire NET_240;
    wire NET_241;
    wire NET_242;
    wire NET_243;
    wire NET_244;
    wire NET_245;
    wire NET_246;
    wire NET_247;
    wire NET_248;
    wire NET_249;
    wire NET_250;
    wire NET_252;
    wire NET_253;
    wire NET_254;
    wire NET_255;
    wire NET_256;
    wire NET_257;
    wire NET_258;
    wire NET_259;
    wire NET_260;
    wire NET_261;
    wire NET_262;
    wire NET_263;
    wire NET_264;
    wire NET_266;
    wire NET_267;
    wire NET_268;
    wire NET_269;
    wire NET_270;
    wire NET_271;
    wire NET_272;
    wire NET_273;
    wire NET_274;
    wire NET_275;
    wire NET_276;
    wire NET_277;
    wire NET_278;
    wire NET_279;
    wire NET_280;
    wire NET_281;
    wire NET_282;
    wire NET_283;
    wire NET_284;
    wire NET_285;
    wire NET_286;
    wire NET_287;
    wire NET_288;
    wire NET_289;
    wire NET_290;
    wire NET_291;
    wire NET_292;
    wire NET_293;
    wire NET_296;
    wire NET_297;
    wire NET_298;
    wire NET_299;
    wire NET_300;
    wire NET_301;
    wire NET_302;
    wire NET_303;
    wire NET_304;
    wire NET_305;
    wire NET_306;
    wire NET_307;
    wire NET_308;
    wire NET_309;
    wire NET_310;
    wire NET_311;
    wire NET_312;
    wire NET_313;
    wire NET_314;
    wire NET_315;
    wire NET_316;
    wire NET_317;
    wire NET_318;
    wire NET_319;
    wire NET_320;
    wire NET_321;
    wire NET_322;
    wire NET_323;
    wire NET_324;
    wire NET_325;
    wire NET_326;
    wire NET_327;
    wire NET_328;
    wire NET_329;
    wire NET_330;
    wire NET_331;
    wire NET_332;
    wire NET_333;
    wire NET_334;
    wire NET_335;
    wire NET_336;
    wire NET_337;
    input wire PCDU;
    input wire PHS4_n;
    input wire PINC;
    input wire PRINC;
    input wire PTWOX;
    input wire R15;
    input wire R6;
    input wire RADRG;
    input wire RADRZ;
    input wire RAND0;
    input wire RBSQ;
    input wire RRPA;
    input wire RUPT0;
    input wire RUPT1;
    input wire SHIFT;
    output wire ST1;
    output wire ST2;
    inout wire ST2_n;
    input wire STBE;
    input wire STBF;
    input wire STFET1_n;
    input wire SU0;
    input wire T01;
    input wire T01_n;
    input wire T02;
    input wire T02_n;
    input wire T03;
    input wire T03_n;
    input wire T04;
    input wire T04_n;
    input wire T05;
    input wire T06;
    input wire T06_n;
    input wire T07;
    input wire T07_n;
    input wire T08;
    input wire T08_n;
    input wire T09;
    input wire T10;
    input wire T10_n;
    input wire T11;
    input wire T11_n;
    input wire T12;
    input wire T12USE_n;
    input wire TL15;
    output wire TSGU_n;
    input wire VCC;
    input wire WAND0;
    wire __A06_1__A2X_n;
    wire __A06_1__BXVX;
    wire __A06_1__CGMC;
    wire __A06_1__CLXC;
    wire __A06_1__DVXP1;
    wire __A06_1__L2GD_n;
    wire __A06_1__MCRO_n;
    wire __A06_1__MONEX;
    wire __A06_1__PIFL_n;
    wire __A06_1__RB1F;
    wire __A06_1__RB_n;
    wire __A06_1__RCH_n;
    wire __A06_1__RC_n;
    wire __A06_1__RG_n;
    wire __A06_1__RU_n;
    wire __A06_1__TOV_n;
    wire __A06_1__TWOX;
    wire __A06_1__WB_n;
    wire __A06_1__WG_n;
    wire __A06_1__WQ_n;
    wire __A06_1__WSC_n;
    wire __A06_1__WYD_n;
    wire __A06_1__WY_n;
    wire __A06_1__WZ_n;
    wire __A06_1__ZAP;
    wire __A06_1__ZAP_n;
    wire __A06_1__ZIP;
    wire __A06_1__ZIPCI;
    wire __A06_2__10XP15;
    wire __A06_2__10XP9;
    wire __A06_2__6XP10;
    wire __A06_2__6XP12;
    wire __A06_2__7XP10;
    wire __A06_2__7XP11;
    wire __A06_2__7XP15;
    wire __A06_2__7XP7;
    wire __A06_2__8XP4;
    wire __A06_2__CI_n;
    wire __A06_2__MOUT;
    wire __A06_2__NEAC;
    wire __A06_2__PONEX;
    wire __A06_2__POUT;
    wire __A06_2__PSEUDO;
    wire __A06_2__R1C_n;
    wire __A06_2__RB1_n;
    wire __A06_2__RB_n;
    wire __A06_2__RC_n;
    wire __A06_2__RDBANK;
    wire __A06_2__RPTSET;
    wire __A06_2__RUS_n;
    wire __A06_2__RU_n;
    wire __A06_2__RZ_n;
    wire __A06_2__WA_n;
    wire __A06_2__WG_n;
    wire __A06_2__WOVR;
    wire __A06_2__WSC_n;
    wire __A06_2__WS_n;
    wire __A06_2__ZOUT;
    input wire n10XP1;
    input wire n10XP8;
    input wire n11XP2;
    input wire n1XP10;
    input wire n2XP3;
    input wire n2XP5;
    input wire n2XP7;
    input wire n2XP8;
    input wire n3XP2;
    input wire n3XP6;
    input wire n3XP7;
    input wire n4XP11;
    input wire n5XP12;
    input wire n5XP15;
    input wire n5XP21;
    input wire n5XP28;
    input wire n5XP4;
    input wire n6XP5;
    input wire n6XP8;
    output wire n7XP14;
    input wire n7XP19;
    input wire n7XP4;
    input wire n7XP9;
    inout wire n8PP4;
    input wire n8XP6;
    input wire n9XP1;
    input wire n9XP5;

    pullup R6001(NET_282);
    pullup R6002(__A06_1__A2X_n);
    pullup R6003(__A06_1__RB_n);
    pullup R6004(__A06_1__WYD_n);
    pullup R6005(NET_268);
    pullup R6006(__A06_1__WYD_n);
    pullup R6007(__A06_1__RG_n);
    pullup R6008(__A06_1__WB_n);
    pullup R6009(__A06_1__RU_n);
    pullup R6010(__A06_1__WZ_n);
    pullup R6011(__A06_1__TOV_n);
    pullup R6012(__A06_1__WSC_n);
    pullup R6013(__A06_1__WG_n);
    pullup R6014(NET_259);
    pullup R6015(NET_223);
    pullup R6016(MONEX_n);
    pullup R6017(__A06_2__RB1_n);
    pullup R6018(__A06_2__R1C_n);
    pullup R6019(n8PP4);
    pullup R6020(NET_203);
    pullup R6021(__A06_2__WS_n);
    pullup R6022(NET_208);
    pullup R6023(__A06_2__CI_n);
    pullup R6024(__A06_2__WA_n);
    pullup R6025(NET_240);
    pullup R6026(ST2_n);
    pullup R6027(__A06_2__RZ_n);
    pullup R6028(__A06_1__RC_n);
    U74HC27 U6001(T04, T07, NET_285, NET_286, NET_287, NET_301, GND, NET_300, T01, T03, T05, NET_284, T10, VCC, SIM_RST);
    U74HC02 U6002(NET_285, NET_284, DV376_n, NET_286, T01_n, DV1376_n, GND, T04_n, DV4_n, NET_287, MP1_n, NET_282, NET_283, VCC, SIM_RST);
    U74HC27 U6003(T07, T09, L15A_n, L02A_n, L01_n, NET_299, GND, NET_315, T05, T08, T11, NET_298, T11, VCC, SIM_RST);
    U74LVC07 U6004(NET_300, NET_282, NET_298, NET_282, NET_309, __A06_1__A2X_n, GND, __A06_1__RB_n, NET_308, __A06_1__WYD_n, NET_310, __A06_1__WY_n, NET_305, VCC, SIM_RST);
    U74HC02 U6005(NET_334, NET_283, n2XP7, __A06_1__L2GD_n, __A06_1__ZIP, __A06_1__DVXP1, GND, __A06_1__DVXP1, NET_303, NET_310, NET_306, NET_302, NET_304, VCC, SIM_RST);
    U74HC04 U6006(L01_n, NET_297, L02A_n, NET_330, L15A_n, NET_335, GND, __A06_1__DVXP1, NET_301, __A06_1__ZIP, NET_334, NET_332, NET_331, VCC, SIM_RST);
    U74HC27 U6007(n7XP19, __A06_1__ZIP, __A06_1__DVXP1, NET_273, RBSQ, NET_308, GND, NET_311, NET_297, NET_330, NET_335, NET_309, __A06_1__DVXP1, VCC, SIM_RST);
    U74HC27 U6008(NET_335, NET_297, NET_334, NET_302, NET_306, NET_305, GND, NET_331, NET_306, NET_302, L02A_n, NET_302, L02A_n, VCC, SIM_RST);
    U74HC02 U6009(NET_303, NET_334, NET_304, NET_307, NET_334, NET_332, GND, NET_315, DV376_n, NET_272, DV1376_n, T02_n, NET_333, VCC, SIM_RST);
    U74HC04 U6010(NET_307, __A06_1__MCRO_n, NET_277, NET_292, NET_275, NET_296, GND, __A06_1__ZAP, __A06_1__ZAP_n, NET_317, NET_315, __A06_1__MONEX, MONEX_n, VCC, SIM_RST);
    U74HC27 U6011(NET_334, NET_332, NET_331, NET_311, NET_334, NET_273, GND, NET_306, NET_330, L15A_n, L01_n, __A06_1__ZIPCI, NET_299, VCC, SIM_RST);
    U74HC02 U6012(NET_277, NET_272, NET_333, NET_275, NET_274, DIVSTG, GND, T08, T10, NET_266, MP1_n, NET_268, NET_271, VCC, SIM_RST);
    U74HC27 U6013(T06, T09, DV376_n, NET_276, T12USE_n, NET_274, GND, NET_267, T02, T04, T06, NET_276, T12, VCC, SIM_RST);
    U74LVC07 U6014(NET_267, NET_268, NET_266, NET_268, NET_291, __A06_1__WYD_n, GND, __A06_1__RG_n, NET_288, __A06_1__WB_n, NET_293, __A06_1__RU_n, NET_281, VCC, SIM_RST);
    U74HC02 U6015(NET_270, T01, T03, NET_269, NET_270, MP3_n, GND, NET_271, NET_269, __A06_1__ZAP_n, n5XP28, NET_292, TSGU_n, VCC, SIM_RST);
    U74HC02 U6016(NET_291, NET_292, n5XP12, NET_278, RRPA, n5XP4, GND, n5XP15, n3XP6, __A06_1__WQ_n, n9XP5, n6XP8, NET_337, VCC, SIM_RST);
    U74HC4002 U6017(NET_288, n5XP4, RADRG, NET_292, n5XP28, NET_289, GND, NET_290, n5XP28, n1XP10, NET_296, n2XP3, NET_293, VCC, SIM_RST);
    U74HC4002 U6018(NET_281, NET_296, __A06_1__ZAP, n5XP12, n6XP5, NET_279, GND, NET_280, PRINC, DINC_n, MINC, DINC, NET_231, VCC, SIM_RST);
    U74LVC07 U6019(NET_278, __A06_1__WZ_n, NET_336, __A06_1__TOV_n, NET_337, __A06_1__WSC_n, GND, __A06_1__WG_n, NET_316, NET_259, NET_264, NET_259, NET_263, VCC, SIM_RST);
    U74HC27 U6020(n6XP5, n3XP2, BR1_n, PHS4_n, TSGU_n, __A06_1__RB1F, GND, __A06_1__CLXC, TSGU_n, BR1, PHS4_n, NET_336, n9XP5, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U6021(NET_316, n6XP8, n6XP8, __A06_1__PIFL_n, __A06_1__DVXP1, NET_312, GND, PTWOX, __A06_1__MONEX, NET_314, __A06_1__MONEX, B15X, NET_313, VCC, SIM_RST);
    U74HC27 U6022(__A06_1__PIFL_n, NET_317, STBE, n1XP10, STBF, NET_319, GND, NET_264, NET_261, NET_260, INCR0, NET_312, T02, VCC, SIM_RST);
    U74HC04 U6023(NET_314, __A06_1__TWOX, NET_313, __A06_1__BXVX, NET_327, NET_328, GND, NET_329, NET_328, NET_326, NET_329, NET_323, NET_326, VCC, SIM_RST);
    U74HC02 U6024(__A06_1__CGMC, NET_319, NET_327, NET_325, __A06_1__CGMC, NET_318, GND, NET_325, NET_319, NET_327, BR1, AUG0_n, NET_261, VCC, SIM_RST);
    U74HC04 U6025(NET_323, NET_322, NET_322, NET_320, NET_320, NET_321, GND, NET_318, NET_321, NET_224, NET_222, NET_233, __A06_2__7XP10, VCC, SIM_RST);
    U74HC02 U6026(NET_260, DIM0_n, BR12B_n, NET_263, PINC, NET_262, GND, BR12B_n, DINC_n, NET_262, T06_n, NET_259, __A06_2__6XP10, VCC, SIM_RST);
    U74HC02 U6027(NET_218, MINC, MCDU, NET_216, AUG0_n, BR1_n, GND, DIM0_n, BR1B2B_n, NET_215, BR1B2B_n, DINC_n, NET_217, VCC, SIM_RST);
    U74HC27 U6028(NET_216, NET_215, BR1B2B_n, CDUSTB_n, DINC_n, __A06_2__POUT, GND, __A06_2__MOUT, BR12B_n, CDUSTB_n, DINC_n, NET_219, NET_217, VCC, SIM_RST);
    U74LVC07 U6029(NET_218, NET_223, NET_219, NET_223, NET_224, MONEX_n, GND, __A06_2__WA_n, NET_213, __A06_2__RB1_n, NET_233, __A06_2__R1C_n, NET_236, VCC, SIM_RST);
    U74HC02 U6030(NET_222, T06_n, NET_223, NET_220, PCDU, MCDU, GND, T06_n, NET_220, __A06_2__6XP12, NET_209, T07_n, NET_212, VCC, SIM_RST);
    U74HC27 U6031(BR2_n, DINC_n, DAS0, DAS1, MSU0, NET_209, GND, NET_213, NET_212, __A06_2__7XP7, NET_207, __A06_2__ZOUT, CDUSTB_n, VCC, SIM_RST);
    U74HC02 U6032(NET_214, DV4_n, BR1B2B, __A06_2__7XP7, T07_n, NET_210, GND, WAND0, INOTLD, NET_235, T07_n, NET_235, n7XP14, VCC, SIM_RST);
    U74HC27 U6033(NET_214, WAND0, DAS1_n, T07_n, BR1B2_n, __A06_2__7XP10, GND, __A06_2__7XP11, DAS1_n, T07_n, BR12B_n, NET_210, RAND0, VCC, SIM_RST);
    U74HC04 U6034(__A06_2__7XP11, NET_236, NET_194, __A06_2__PONEX, ST2_n, ST2, GND, ST1, NET_249, NET_246, __A06_2__PSEUDO, NET_247, __A06_2__RDBANK, VCC, SIM_RST);
    U74HC02 U6035(__A06_2__7XP15, NET_227, T07_n, NET_230, NET_231, T07_n, GND, PRINC, INKL, NET_229, IC9, DXCH0, NET_191, VCC, SIM_RST);
    U74HC27 U6036(PCDU, MCDU, n7XP9, n11XP2, __A06_2__7XP15, __A06_2__RUS_n, GND, NET_232, NET_230, NET_238, NET_207, NET_227, SHIFT, VCC, SIM_RST);
    U74LVC07 U6037(NET_232, __A06_2__RU_n, NET_187, __A06_2__WSC_n, NET_188, __A06_2__WG_n, GND, __A06_2__RB_n, NET_190, n8PP4, NET_183, n8PP4, NET_181, VCC, SIM_RST);
    U74HC27 U6038(NET_229, T07_n, T04_n, MON_n, FETCH1, NET_189, GND, NET_187, __A06_2__WOVR, NET_189, NET_244, __A06_2__WOVR, MONPCH, VCC, SIM_RST);
    U74HC02 U6039(NET_188, __A06_2__WOVR, NET_244, NET_244, T07_n, NET_191, GND, __A06_2__10XP9, NET_244, NET_190, T08_n, n8PP4, __A06_2__8XP4, VCC, SIM_RST);
    U74HC27 U6040(RUPT1, DAS1, IC17, MASK0, IC11, NET_181, GND, NET_182, IC6, IC7, DV4B1B, NET_183, DV4_n, VCC, SIM_RST);
    U74LVC07 U6041(NET_182, n8PP4, NET_185, NET_203, NET_184, NET_203, GND, __A06_2__WS_n, NET_204, NET_208, NET_202, NET_208, NET_205, VCC, SIM_RST);
    U74HC27 U6042(T08_n, RUPT0, NET_203, R6, R15, NET_204, GND, NET_205, ADS0, IC11, NET_206, NET_185, DAS0, VCC, SIM_RST);
    U74HC02 U6043(NET_184, MP1, DV1376, NET_201, MP3_n, BR1_n, GND, NET_201, CCS0, NET_202, T11_n, NET_208, NET_207, VCC, SIM_RST);
    U74HC02 U6044(NET_206, DAS1_n, BR2_n, NET_193, __A06_1__ZIPCI, __A06_2__6XP12, GND, CCS0_n, BR1B2B_n, NET_199, T10_n, NDXX1_n, EXT, VCC, SIM_RST);
    U74HC27 U6045(T03_n, DAS1_n, NET_243, NET_238, n2XP5, NET_257, GND, NET_252, IC7, DCS0, SU0, NET_238, ADS0, VCC, SIM_RST);
    U74HC4002 U6046(NET_194, n8XP6, n7XP4, n10XP8, __A06_2__6XP10, NET_195, GND, NET_196, IC6, DCA0, AD0, NET_199, NET_200, VCC, SIM_RST);
    U74LVC07 U6047(NET_193, __A06_2__CI_n, NET_257, __A06_2__WA_n, NET_258, __A06_2__RC_n, GND, NET_240, NET_252, NET_240, NET_253, ST2_n, NET_256, VCC, SIM_RST);
    U74HC02 U6048(__A06_2__10XP9, T10_n, NET_200, NET_242, IC6, IC7, GND, T10_n, NET_242, NET_243, T10_n, NET_240, NET_239, VCC, SIM_RST);
    U74HC02 U6049(NET_258, NET_239, __A06_2__7XP7, NET_253, NET_241, DV4B1B, GND, CCS0_n, BR12B_n, NET_241, T10_n, MP1_n, __A06_2__10XP15, VCC, SIM_RST);
    U74HC27 U6050(__A06_2__8XP4, __A06_2__10XP15, __A06_2__8XP4, RADRZ, n9XP1, NET_248, GND, __A06_2__NEAC, NET_250, TL15, GOJAM, NET_256, RADRZ, VCC, SIM_RST);
    wire U6051_9_NC;
    wire U6051_10_NC;
    wire U6051_11_NC;
    wire U6051_12_NC;
    wire U6051_13_NC;
    U74HC4002 U6051(NET_249, n2XP8, n10XP1, MP0T10, __A06_2__10XP15, NET_254, GND, NET_255, U6051_9_NC, U6051_10_NC, U6051_11_NC, U6051_12_NC, U6051_13_NC, VCC, SIM_RST);
    wire U6052_10_NC;
    wire U6052_11_NC;
    wire U6052_12_NC;
    wire U6052_13_NC;
    U74LVC07 U6052(NET_248, __A06_2__RZ_n, NET_246, __A06_2__RPTSET, NET_247, __A06_2__RU_n, GND, __A06_1__RC_n, NET_324, U6052_10_NC, U6052_11_NC, U6052_12_NC, U6052_13_NC, VCC, SIM_RST);
    U74HC02 #(1, 0, 0, 0) U6053(NET_250, MP0T10, __A06_2__NEAC, NET_245, RADRZ, __A06_2__PSEUDO, GND, T06_n, STFET1_n, __A06_2__RDBANK, __A06_1__ZIPCI, n3XP7, NET_324, VCC, SIM_RST);
    wire U6054_8_NC;
    wire U6054_9_NC;
    wire U6054_10_NC;
    wire U6054_11_NC;
    U74HC27 #(1, 0, 0) U6054(NET_245, GOJAM, n3XP7, n5XP21, n4XP11, __A06_1__RCH_n, GND, U6054_8_NC, U6054_9_NC, U6054_10_NC, U6054_11_NC, __A06_2__PSEUDO, RADRG, VCC, SIM_RST);
endmodule