`timescale 1ns/1ps
`default_nettype none

module fixed_erasable_memory(VCC, GND, SIM_RST, SIM_CLK, ROPER, ROPES, ROPET, HIMOD, LOMOD, STR14, STR58, STR912, STR19, STR210, STR311, STR412, SETAB, SETCD, RESETA, RESETB, RESETC, RESETD, CLROPE, IL07, IL06, IL05, IL04, IL03, IL02, IL01, SBF, XB7E, XB1E, XB2E, XB3E, XB4E, XB5E, XB6E, XT7E, XT1E, XT2E, XT3E, XT4E, XT5E, XT6E, YB3E, YB1E, YB2E, YT7E, YT1E, YT2E, YT3E, YT4E, YT5E, YT6E, GEMP, GEM01, GEM02, GEM03, GEM04, GEM05, GEM06, GEM07, GEM08, GEM09, GEM10, GEM11, GEM12, GEM13, GEM14, GEM16, SETEK, RSTKX_n, RSTKY_n, SBE, REX, REY, WEX, WEY, ZID, SAP, SA01, SA02, SA03, SA04, SA05, SA06, SA07, SA08, SA09, SA10, SA11, SA12, SA13, SA14, SA16);
    input wire VCC;
    input wire GND;
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire CLROPE;
    input wire GEM01;
    input wire GEM02;
    input wire GEM03;
    input wire GEM04;
    input wire GEM05;
    input wire GEM06;
    input wire GEM07;
    input wire GEM08;
    input wire GEM09;
    input wire GEM10;
    input wire GEM11;
    input wire GEM12;
    input wire GEM13;
    input wire GEM14;
    input wire GEM16;
    input wire GEMP;
    input wire HIMOD;
    input wire IL01;
    input wire IL02;
    input wire IL03;
    input wire IL04;
    input wire IL05;
    input wire IL06;
    input wire IL07;
    input wire LOMOD;
    input wire RESETA;
    input wire RESETB;
    input wire RESETC;
    input wire RESETD;
    input wire REX;
    input wire REY;
    input wire ROPER;
    input wire ROPES;
    input wire ROPET;
    input wire RSTKX_n;
    input wire RSTKY_n;
    output wire SA01; //FPGA#wor
    output wire SA02; //FPGA#wor
    output wire SA03; //FPGA#wor
    output wire SA04; //FPGA#wor
    output wire SA05; //FPGA#wor
    output wire SA06; //FPGA#wor
    output wire SA07; //FPGA#wor
    output wire SA08; //FPGA#wor
    output wire SA09; //FPGA#wor
    output wire SA10; //FPGA#wor
    output wire SA11; //FPGA#wor
    output wire SA12; //FPGA#wor
    output wire SA13; //FPGA#wor
    output wire SA14; //FPGA#wor
    output wire SA16; //FPGA#wor
    output wire SAP; //FPGA#wor
    input wire SBE;
    input wire SBF;
    input wire SETAB;
    input wire SETCD;
    input wire SETEK;
    input wire STR14;
    input wire STR19;
    input wire STR210;
    input wire STR311;
    input wire STR412;
    input wire STR58;
    input wire STR912;
    input wire WEX;
    input wire WEY;
    input wire XB1E;
    input wire XB2E;
    input wire XB3E;
    input wire XB4E;
    input wire XB5E;
    input wire XB6E;
    input wire XB7E;
    input wire XT1E;
    input wire XT2E;
    input wire XT3E;
    input wire XT4E;
    input wire XT5E;
    input wire XT6E;
    input wire XT7E;
    input wire YB1E;
    input wire YB2E;
    input wire YB3E;
    input wire YT1E;
    input wire YT2E;
    input wire YT3E;
    input wire YT4E;
    input wire YT5E;
    input wire YT6E;
    input wire YT7E;
    input wire ZID;
    wire __B01_1__CQA;
    wire __B01_1__CQB;
    wire __B01_1__CQC;
    wire __B01_1__FADDR1;
    wire __B01_1__FADDR10;
    wire __B01_1__FADDR11;
    wire __B01_1__FADDR12;
    wire __B01_1__FADDR13;
    wire __B01_1__FADDR14;
    wire __B01_1__FADDR15;
    wire __B01_1__FADDR16;
    wire __B01_1__FADDR2;
    wire __B01_1__FADDR3;
    wire __B01_1__FADDR4;
    wire __B01_1__FADDR5;
    wire __B01_1__FADDR6;
    wire __B01_1__FADDR7;
    wire __B01_1__FADDR8;
    wire __B01_1__FADDR9;
    wire __B01_1__NOROPE;
    wire __B01_1__QUARTERA;
    wire __B01_1__QUARTERB;
    wire __B01_1__QUARTERC;
    wire __B01_2__EDESTROY;
    wire __B01_2__ES01_n;
    wire __B01_2__ES02_n;
    wire __B01_2__ES03_n;
    wire __B01_2__ES04_n;
    wire __B01_2__ES05_n;
    wire __B01_2__ES06_n;
    wire __B01_2__ES07_n;
    wire __B01_2__ES08_n;
    wire __B01_2__ES09_n;
    wire __B01_2__ES10_n;
    wire __B01_2__ES11_n;
    wire __B01_2__RADDR1;
    wire __B01_2__RADDR10;
    wire __B01_2__RADDR11;
    wire __B01_2__RADDR2;
    wire __B01_2__RADDR3;
    wire __B01_2__RADDR4;
    wire __B01_2__RADDR5;
    wire __B01_2__RADDR6;
    wire __B01_2__RADDR7;
    wire __B01_2__RADDR8;
    wire __B01_2__RADDR9;
    wire __B01_2__RESETK;
    wire __B01_NET_100;
    wire __B01_NET_101;
    wire __B01_NET_102;
    wire __B01_NET_103;
    wire __B01_NET_105;
    wire __B01_NET_106;
    wire __B01_NET_107;
    wire __B01_NET_108;
    wire __B01_NET_109;
    wire __B01_NET_110;
    wire __B01_NET_114;
    wire __B01_NET_115;
    wire __B01_NET_116;
    wire __B01_NET_119;
    wire __B01_NET_120;
    wire __B01_NET_121;
    wire __B01_NET_122;
    wire __B01_NET_123;
    wire __B01_NET_124;
    wire __B01_NET_125;
    wire __B01_NET_127;
    wire __B01_NET_128;
    wire __B01_NET_131;
    wire __B01_NET_132;
    wire __B01_NET_133;
    wire __B01_NET_134;
    wire __B01_NET_135;
    wire __B01_NET_136;
    wire __B01_NET_137;
    wire __B01_NET_138;
    wire __B01_NET_139;
    wire __B01_NET_140;
    wire __B01_NET_141;
    wire __B01_NET_142;
    wire __B01_NET_143;
    wire __B01_NET_144;
    wire __B01_NET_146;
    wire __B01_NET_147;
    wire __B01_NET_148;
    wire __B01_NET_149;
    wire __B01_NET_150;
    wire __B01_NET_152;
    wire __B01_NET_158;
    wire __B01_NET_176;
    wire __B01_NET_177;
    wire __B01_NET_178;
    wire __B01_NET_179;
    wire __B01_NET_180;
    wire __B01_NET_181;
    wire __B01_NET_182;
    wire __B01_NET_183;
    wire __B01_NET_186;
    wire __B01_NET_189;
    wire __B01_NET_190;
    wire __B01_NET_191;
    wire __B01_NET_192;
    wire __B01_NET_195;
    wire __B01_NET_196;
    wire __B01_NET_197;
    wire __B01_NET_198;
    wire __B01_NET_199;
    wire __B01_NET_201;
    wire __B01_NET_202;
    wire __B01_NET_204;
    wire __B01_NET_208;
    wire __B01_NET_210;
    wire __B01_NET_212;
    wire __B01_NET_213;
    wire __B01_NET_217;
    wire __B01_NET_218;
    wire __B01_NET_224;
    wire __B01_NET_225;
    wire __B01_NET_226;
    wire __B01_NET_227;
    wire __B01_NET_228;
    wire __B01_NET_229;
    wire __B01_NET_230;
    wire __B01_NET_231;
    wire __B01_NET_232;
    wire __B01_NET_233;
    wire __B01_NET_234;
    wire __B01_NET_235;
    wire __B01_NET_236;
    wire __B01_NET_239;
    wire __B01_NET_240;
    wire __B01_NET_241;
    wire __B01_NET_242;
    wire __B01_NET_243;
    wire __B01_NET_245;
    wire __B01_NET_246;
    wire __B01_NET_247;
    wire __B01_NET_249;
    wire __B01_NET_251;
    wire __B01_NET_253;
    wire __B01_NET_95;
    wire __B01_NET_97;
    wire __B01_NET_98;
    wire __B01_NET_99;

    pulldown R31001(SAP);
    pulldown R31002(SA01);
    pulldown R31003(SA02);
    pulldown R31004(SA03);
    pulldown R31005(SA04);
    pulldown R31006(SA05);
    pulldown R31007(SA06);
    pulldown R31008(SA07);
    pulldown R31009(SA08);
    pulldown R31010(SA09);
    pulldown R31011(SA10);
    pulldown R31012(SA11);
    pulldown R31013(SA12);
    pulldown R31014(SA13);
    pulldown R31015(SA14);
    pulldown R31016(SA16);
    SST39VF200A U31001(__B01_1__FADDR16, __B01_1__FADDR15, __B01_1__FADDR14, __B01_1__FADDR13, __B01_1__FADDR12, __B01_1__FADDR11, __B01_1__FADDR10, __B01_1__FADDR9,  ,  , VCC,  ,  ,  ,  ,  ,  , __B01_1__FADDR8, __B01_1__FADDR7, __B01_1__FADDR6, __B01_1__FADDR5, __B01_1__FADDR4, __B01_1__FADDR3, __B01_1__FADDR2, __B01_1__FADDR1, __B01_NET_158, GND, __B01_NET_110, SAP, SA08, SA01, SA09, SA02, SA10, SA03, SA11, VCC, SA04, SA12, SA05, SA13, SA06, SA14, SA07, SA16, GND,  , GND, SIM_RST, SIM_CLK); //FPGA#inputs:EPCS_DATA;FPGA#outputs:EPCS_CSN,EPCS_DCLK,EPCS_ASDI;FPGA#OD:29,30,31,32,33,34,35,36,38,39,40,41,42,43,44,45
    U74HC04 U31002(ROPER, __B01_NET_176, ROPES, __B01_NET_189, ROPET, __B01_NET_144, GND, __B01_NET_177, STR14, __B01_NET_180, STR58, __B01_NET_143, STR912, VCC, SIM_RST, SIM_CLK);
    U74HC27 U31003(__B01_NET_144, LOMOD, ROPER, __B01_NET_146, __B01_NET_186, __B01_1__FADDR15, GND, __B01_NET_146, ROPES, LOMOD, STR14, __B01_1__FADDR16, STR14, VCC, SIM_RST, SIM_CLK);
    U74HC27 U31004(ROPET, HIMOD, ROPER, LOMOD, STR14, __B01_NET_149, GND, __B01_NET_148, ROPET, LOMOD, __B01_NET_177, __B01_NET_186, STR912, VCC, SIM_RST, SIM_CLK);
    U74HC02 U31005(__B01_NET_150, __B01_NET_189, __B01_NET_143, __B01_NET_147, __B01_NET_176, HIMOD, GND, HIMOD, STR58, __B01_NET_179, LOMOD, __B01_NET_180, __B01_NET_178, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U31006(__B01_1__FADDR14, __B01_NET_150, __B01_NET_149, __B01_NET_148, __B01_NET_147,  , GND,  , __B01_NET_152, __B01_NET_183, __B01_NET_182, __B01_NET_181, __B01_1__FADDR13, VCC, SIM_RST, SIM_CLK);
    U74HC27 U31007(ROPES, HIMOD, ROPES, LOMOD, STR14, __B01_NET_183, GND, __B01_NET_182, __B01_NET_189, HIMOD, __B01_NET_143, __B01_NET_152, STR912, VCC, SIM_RST, SIM_CLK);
    U74HC27 U31008(__B01_NET_189, LOMOD, RSTKX_n, RSTKY_n, ZID, __B01_2__RESETK, GND, __B01_1__NOROPE, ROPER, ROPES, ROPET, __B01_NET_181, __B01_NET_177, VCC, SIM_RST, SIM_CLK);
    U74HC02 U31009(__B01_1__FADDR12, __B01_NET_179, __B01_NET_178, __B01_1__FADDR11, STR210, STR19, GND, STR19, STR311, __B01_1__FADDR10, __B01_1__QUARTERB, __B01_1__QUARTERA, __B01_1__FADDR9, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31010(__B01_1__FADDR8, __B01_1__QUARTERA, __B01_1__QUARTERC, __B01_NET_116, __B01_NET_115, __B01_1__QUARTERA, GND, __B01_NET_116, __B01_1__CQA, __B01_1__QUARTERA, __B01_NET_102, __B01_NET_99, __B01_NET_115, VCC, SIM_RST, SIM_CLK);
    U74HC04 U31011(IL07, __B01_1__FADDR7, IL06, __B01_1__FADDR6, IL05, __B01_1__FADDR5, GND, __B01_1__FADDR4, IL04, __B01_1__FADDR3, IL03, __B01_1__FADDR2, IL02, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1) U31012(IL01, __B01_1__FADDR1, __B01_NET_114, __B01_NET_110, SETAB, __B01_NET_102, GND, __B01_NET_99, RESETB, __B01_NET_225, __B01_NET_224, __B01_NET_98, __B01_NET_101, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U31013(__B01_NET_158, STR19, STR210, STR311, STR412,  , GND,  , XB1E, XB3E, XB5E, XB7E, __B01_2__ES01_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31014(__B01_NET_97, RESETA, __B01_NET_100, __B01_NET_95, __B01_NET_97, __B01_NET_101, GND, __B01_NET_95, RESETA, __B01_NET_101, __B01_NET_102, __B01_NET_137, __B01_NET_136, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1) U31015(__B01_NET_98, __B01_NET_107, __B01_NET_107, __B01_NET_109, __B01_NET_139, __B01_NET_108, GND, __B01_NET_103, __B01_NET_108, __B01_NET_105, __B01_NET_103, __B01_NET_140, __B01_NET_105, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1) U31016(__B01_NET_109, __B01_NET_100, RESETA, __B01_NET_137, SETCD, __B01_NET_142, GND, __B01_NET_135, RESETD, __B01_1__CQA, __B01_NET_141, __B01_NET_218, ZID, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U31017(__B01_NET_106, __B01_NET_136, __B01_1__QUARTERB, __B01_1__QUARTERB, __B01_NET_106, __B01_1__CQB, GND, __B01_NET_133, __B01_1__QUARTERC, __B01_NET_134, __B01_NET_134, __B01_1__CQC, __B01_1__QUARTERC, VCC, SIM_RST, SIM_CLK);
    U74HC02 U31018(__B01_NET_133, __B01_NET_142, __B01_NET_135, __B01_NET_141, CLROPE, __B01_NET_97, GND, YB1E, YB3E, __B01_2__ES07_n, YB2E, YB3E, __B01_2__ES08_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U31019(__B01_2__ES02_n, XB2E, XB3E, XB6E, XB7E,  , GND,  , XB4E, XB5E, XB6E, XB7E, __B01_2__ES03_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U31020(__B01_2__ES04_n, XT1E, XT3E, XT5E, XT7E,  , GND,  , XT2E, XT3E, XT6E, XT7E, __B01_2__ES05_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U31021(__B01_2__ES06_n, XT4E, XT5E, XT6E, XT7E,  , GND,  , YT1E, YT3E, YT5E, YT7E, __B01_2__ES09_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U31022(__B01_2__ES10_n, YT2E, YT3E, YT6E, YT7E,  , GND,  , YT4E, YT5E, YT6E, YT7E, __B01_2__ES11_n, VCC, SIM_RST, SIM_CLK);
    U74HC244 U31023(__B01_NET_218, GEMP, SA07, GEM01, SA06, GEM02, SA05, GEM03, SA04, GND, GEM04, SA03, GEM05, SA02, GEM06, SA01, GEM07, SAP, __B01_NET_218, VCC, SIM_RST, SIM_CLK); //FPGA#OD:3,5,7,9,12,14,16,18
    U74HC244 U31024(__B01_NET_218, GEM08, SA16, GEM09, SA14, GEM10, SA13, GEM11, SA12, GND, GEM12, SA11, GEM13, SA10, GEM14, SA09, GEM16, SA08, __B01_NET_218, VCC, SIM_RST, SIM_CLK); //FPGA#OD:3,5,7,9,12,14,16,18
    MR0A16A U31025(__B01_2__RADDR1, __B01_2__RADDR2, __B01_2__RADDR3, __B01_2__RADDR4, __B01_2__RADDR5, GND, SAP, SA01, SA02, SA03, VCC, GND, SA04, SA05, SA06, SA07, __B01_NET_196, __B01_2__RADDR6, __B01_2__RADDR7, __B01_2__RADDR8, __B01_2__RADDR9, __B01_2__RADDR10, __B01_2__RADDR11, GND, GND, GND, VCC,  , SA08, SA09, SA10, SA11, VCC, GND, SA12, SA13, SA14, SA16, GND, GND, __B01_NET_191, GND, GND, GND, SIM_RST, SIM_CLK); //FPGA#bidir:7,8,9,10,13,14,15,16,29,30,31,32,35,36,37,38;FPGA#OD:7,8,9,10,13,14,15,16,29,30,31,32,35,36,37,38
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31026(__B01_NET_234, __B01_NET_195, __B01_NET_192, __B01_NET_197, __B01_2__ES01_n, __B01_NET_253, GND, __B01_NET_197, __B01_2__RADDR1, __B01_NET_190, __B01_NET_190, __B01_2__RESETK, __B01_2__RADDR1, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1) U31027(WEX, __B01_NET_195, WEY, __B01_NET_192, __B01_NET_232, __B01_NET_233, GND, __B01_NET_191, SBE, __B01_NET_253, SETEK, __B01_NET_231, __B01_NET_230, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31028(__B01_NET_201, __B01_2__ES02_n, __B01_NET_253, __B01_NET_202, __B01_NET_201, __B01_2__RADDR2, GND, __B01_NET_202, __B01_2__RESETK, __B01_2__RADDR2, __B01_2__ES03_n, __B01_NET_253, __B01_NET_198, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U31029(__B01_NET_199, __B01_NET_198, __B01_2__RADDR3, __B01_2__RADDR3, __B01_NET_199, __B01_2__RESETK, GND, __B01_2__ES04_n, __B01_NET_253, __B01_NET_246, __B01_NET_246, __B01_2__RADDR4, __B01_NET_247, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31030(__B01_2__RADDR4, __B01_NET_247, __B01_2__RESETK, __B01_NET_245, __B01_2__ES05_n, __B01_NET_253, GND, __B01_NET_245, __B01_2__RADDR5, __B01_NET_243, __B01_NET_243, __B01_2__RESETK, __B01_2__RADDR5, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31031(__B01_NET_251, __B01_2__ES06_n, __B01_NET_253, __B01_NET_249, __B01_NET_251, __B01_2__RADDR6, GND, __B01_NET_249, __B01_2__RESETK, __B01_2__RADDR6, __B01_2__ES07_n, __B01_NET_253, __B01_NET_241, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U31032(__B01_NET_242, __B01_NET_241, __B01_2__RADDR7, __B01_2__RADDR7, __B01_NET_242, __B01_2__RESETK, GND, __B01_2__ES08_n, __B01_NET_253, __B01_NET_239, __B01_NET_239, __B01_2__RADDR8, __B01_NET_240, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31033(__B01_2__RADDR8, __B01_NET_240, __B01_2__RESETK, __B01_NET_212, __B01_2__ES09_n, __B01_NET_253, GND, __B01_NET_212, __B01_2__RADDR9, __B01_NET_210, __B01_NET_210, __B01_2__RESETK, __B01_2__RADDR9, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31034(__B01_NET_217, __B01_2__ES10_n, __B01_NET_253, __B01_NET_213, __B01_NET_217, __B01_2__RADDR10, GND, __B01_NET_213, __B01_2__RESETK, __B01_2__RADDR10, __B01_2__ES11_n, __B01_NET_253, __B01_NET_204, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U31035(__B01_NET_208, __B01_NET_204, __B01_2__RADDR11, __B01_NET_125, CLROPE, __B01_NET_127, GND, __B01_NET_233, __B01_NET_236, __B01_2__EDESTROY, __B01_2__EDESTROY, __B01_NET_230, __B01_NET_229, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31036(__B01_NET_230, __B01_NET_229, __B01_NET_233, __B01_NET_127, RESETB, __B01_NET_140, GND, __B01_NET_127, __B01_NET_139, __B01_NET_138, __B01_NET_138, RESETB, __B01_NET_139, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1) U31037(__B01_NET_231, __B01_NET_224, __B01_NET_125, __B01_1__CQB, __B01_NET_225, __B01_NET_228, GND, __B01_NET_226, __B01_NET_228, __B01_NET_227, __B01_NET_226, __B01_NET_235, __B01_NET_227, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1) U31038(__B01_NET_235, __B01_NET_236, __B01_NET_132, __B01_1__CQC, __B01_NET_124, __B01_NET_128, GND, __B01_NET_119, __B01_NET_128, __B01_NET_121, __B01_NET_119, __B01_NET_120, __B01_NET_121, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31039(__B01_NET_132, CLROPE, __B01_NET_123, __B01_NET_123, RESETC, __B01_NET_120, GND, __B01_NET_123, __B01_NET_124, __B01_NET_122, __B01_NET_122, RESETC, __B01_NET_124, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U31040(__B01_2__RADDR11, __B01_NET_208, __B01_2__RESETK, __B01_NET_232, REX, REY, GND, __B01_NET_234, __B01_2__EDESTROY, __B01_NET_196, __B01_NET_131, __B01_1__NOROPE, __B01_NET_114, VCC, SIM_RST, SIM_CLK);
    U74HC04 U31041(SBF, __B01_NET_131,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
endmodule