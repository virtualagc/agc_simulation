`timescale 1ns/1ps

module crosspoint_ii(VCC, GND, SIM_RST, GOJAM, T01, T01_n, T02, T02_n, T03, T03_n, T04, T04_n, T05, T06, T06_n, T07, T07_n, T08, T08_n, T09, T10, T10_n, T11, T11_n, T12, T12USE_n, PHS4_n, ST2_n, BR1, BR1_n, BR2_n, BR1B2_n, BR12B_n, BR1B2B, BR1B2B_n, INKL, AD0, ADS0, AUG0_n, CCS0, CCS0_n, CDUSTB_n, DAS0, DAS1, DAS1_n, DCA0, DCS0, DIM0_n, DINC, DINC_n, DV1376, DV1376_n, DV376_n, DV4_n, DV4B1B, DXCH0, FETCH1, INCR0, INOTLD, MASK0, MCDU, MINC, MP0T10, MP1, MP1_n, MP3_n, MSU0, NDXX1_n, PCDU, PINC, PRINC, RAND0, RUPT0, RUPT1, SHIFT, STFET1_n, SU0, WAND0, IC6, IC7, IC9, IC11, IC17, B15X, DIVSTG, PTWOX, R6, R15, RADRG, RADRZ, RBSQ, RRPA, STBE, STBF, TL15, L01_n, L02A_n, L15A_n, MON_n, MONPCH, n8PP4, n1XP10, n2XP3, n2XP5, n2XP7, n2XP8, n3XP2, n3XP6, n3XP7, n4XP11, n5XP4, n5XP12, n5XP15, n5XP21, n5XP28, n6XP5, n6XP8, n7XP4, n7XP9, n7XP19, n8XP6, n9XP1, n9XP5, n10XP1, n10XP8, n11XP2, A2X_n, CGMC, CI_n, EXT, L2GD_n, MONEX_n, NEAC, PIFL_n, RB_n, RC_n, RCH_n, RG_n, RU_n, RUS_n, RZ_n, ST1, ST2, TOV_n, TSGU_n, WA_n, WB_n, WG_n, WL_n, WQ_n, WS_n, WSC_n, WY_n, WYD_n, WZ_n, ZAP_n, RPTSET, n7XP14);
    input wire SIM_RST;
    inout wire A2X_n;
    input wire AD0;
    input wire ADS0;
    input wire AUG0_n;
    input wire B15X;
    input wire BR1;
    input wire BR12B_n;
    input wire BR1B2B;
    input wire BR1B2B_n;
    input wire BR1B2_n;
    input wire BR1_n;
    input wire BR2_n;
    input wire CCS0;
    input wire CCS0_n;
    input wire CDUSTB_n;
    output wire CGMC;
    inout wire CI_n;
    input wire DAS0;
    input wire DAS1;
    input wire DAS1_n;
    input wire DCA0;
    input wire DCS0;
    input wire DIM0_n;
    input wire DINC;
    input wire DINC_n;
    input wire DIVSTG;
    input wire DV1376;
    input wire DV1376_n;
    input wire DV376_n;
    input wire DV4B1B;
    input wire DV4_n;
    input wire DXCH0;
    output wire EXT;
    input wire FETCH1;
    input wire GND;
    input wire GOJAM;
    input wire IC11;
    input wire IC17;
    input wire IC6;
    input wire IC7;
    input wire IC9;
    input wire INCR0;
    input wire INKL;
    input wire INOTLD;
    input wire L01_n;
    input wire L02A_n;
    input wire L15A_n;
    output wire L2GD_n;
    input wire MASK0;
    input wire MCDU;
    input wire MINC;
    inout wire MONEX_n;
    input wire MONPCH;
    input wire MON_n;
    input wire MP0T10;
    input wire MP1;
    input wire MP1_n;
    input wire MP3_n;
    input wire MSU0;
    input wire NDXX1_n;
    output wire NEAC;
    wire NET_177;
    wire NET_178;
    wire NET_179;
    wire NET_180;
    wire NET_181;
    wire NET_183;
    wire NET_184;
    wire NET_185;
    wire NET_186;
    wire NET_187;
    wire NET_189;
    wire NET_190;
    wire NET_191;
    wire NET_192;
    wire NET_195;
    wire NET_196;
    wire NET_197;
    wire NET_198;
    wire NET_199;
    wire NET_200;
    wire NET_201;
    wire NET_202;
    wire NET_203;
    wire NET_204;
    wire NET_205;
    wire NET_206;
    wire NET_208;
    wire NET_209;
    wire NET_210;
    wire NET_211;
    wire NET_212;
    wire NET_213;
    wire NET_214;
    wire NET_215;
    wire NET_216;
    wire NET_218;
    wire NET_219;
    wire NET_220;
    wire NET_223;
    wire NET_225;
    wire NET_226;
    wire NET_227;
    wire NET_228;
    wire NET_229;
    wire NET_231;
    wire NET_232;
    wire NET_234;
    wire NET_235;
    wire NET_236;
    wire NET_237;
    wire NET_238;
    wire NET_239;
    wire NET_240;
    wire NET_241;
    wire NET_242;
    wire NET_243;
    wire NET_244;
    wire NET_245;
    wire NET_246;
    wire NET_248;
    wire NET_249;
    wire NET_250;
    wire NET_251;
    wire NET_252;
    wire NET_253;
    wire NET_254;
    wire NET_255;
    wire NET_256;
    wire NET_257;
    wire NET_258;
    wire NET_259;
    wire NET_260;
    wire NET_262;
    wire NET_263;
    wire NET_264;
    wire NET_265;
    wire NET_266;
    wire NET_267;
    wire NET_268;
    wire NET_269;
    wire NET_270;
    wire NET_271;
    wire NET_272;
    wire NET_273;
    wire NET_274;
    wire NET_275;
    wire NET_276;
    wire NET_277;
    wire NET_278;
    wire NET_279;
    wire NET_280;
    wire NET_281;
    wire NET_282;
    wire NET_283;
    wire NET_284;
    wire NET_285;
    wire NET_286;
    wire NET_287;
    wire NET_288;
    wire NET_289;
    wire NET_292;
    wire NET_293;
    wire NET_294;
    wire NET_295;
    wire NET_296;
    wire NET_297;
    wire NET_298;
    wire NET_299;
    wire NET_300;
    wire NET_301;
    wire NET_302;
    wire NET_303;
    wire NET_304;
    wire NET_305;
    wire NET_306;
    wire NET_307;
    wire NET_308;
    wire NET_309;
    wire NET_310;
    wire NET_311;
    wire NET_312;
    wire NET_313;
    wire NET_314;
    wire NET_315;
    wire NET_316;
    wire NET_317;
    wire NET_318;
    wire NET_319;
    wire NET_320;
    wire NET_321;
    wire NET_322;
    wire NET_323;
    wire NET_324;
    wire NET_325;
    wire NET_326;
    wire NET_327;
    wire NET_328;
    wire NET_329;
    wire NET_330;
    wire NET_331;
    wire NET_332;
    wire NET_333;
    input wire PCDU;
    input wire PHS4_n;
    output wire PIFL_n;
    input wire PINC;
    input wire PRINC;
    input wire PTWOX;
    input wire R15;
    input wire R6;
    input wire RADRG;
    input wire RADRZ;
    input wire RAND0;
    input wire RBSQ;
    inout wire RB_n;
    output wire RCH_n;
    inout wire RC_n;
    inout wire RG_n;
    inout wire RPTSET;
    input wire RRPA;
    input wire RUPT0;
    input wire RUPT1;
    output wire RUS_n;
    inout wire RU_n;
    inout wire RZ_n;
    input wire SHIFT;
    output wire ST1;
    output wire ST2;
    inout wire ST2_n;
    input wire STBE;
    input wire STBF;
    input wire STFET1_n;
    input wire SU0;
    input wire T01;
    input wire T01_n;
    input wire T02;
    input wire T02_n;
    input wire T03;
    input wire T03_n;
    input wire T04;
    input wire T04_n;
    input wire T05;
    input wire T06;
    input wire T06_n;
    input wire T07;
    input wire T07_n;
    input wire T08;
    input wire T08_n;
    input wire T09;
    input wire T10;
    input wire T10_n;
    input wire T11;
    input wire T11_n;
    input wire T12;
    input wire T12USE_n;
    input wire TL15;
    inout wire TOV_n;
    output wire TSGU_n;
    input wire VCC;
    input wire WAND0;
    inout wire WA_n;
    inout wire WB_n;
    inout wire WG_n;
    inout wire WL_n;
    output wire WQ_n;
    inout wire WSC_n;
    inout wire WS_n;
    inout wire WYD_n;
    inout wire WY_n;
    inout wire WZ_n;
    output wire ZAP_n;
    wire __A06_1__BXVX;
    wire __A06_1__CGMC;
    wire __A06_1__CLXC;
    wire __A06_1__MCRO_n;
    wire __A06_1__MONEX;
    wire __A06_1__RB1F;
    wire __A06_1__TWOX;
    wire __A06_1__ZAP;
    wire __A06_1__ZIP;
    wire __A06_1__ZIPCI;
    wire __A06_2__10XP15;
    wire __A06_2__10XP9;
    wire __A06_2__6XP10;
    wire __A06_2__6XP12;
    wire __A06_2__7XP10;
    wire __A06_2__7XP11;
    wire __A06_2__7XP15;
    wire __A06_2__7XP7;
    wire __A06_2__8XP4;
    wire __A06_2__MOUT;
    wire __A06_2__PONEX;
    wire __A06_2__POUT;
    wire __A06_2__PSEUDO;
    wire __A06_2__R1C_n;
    wire __A06_2__RB1_n;
    wire __A06_2__RDBANK;
    wire __A06_2__WOVR;
    wire __A06_2__ZOUT;
    input wire n10XP1;
    input wire n10XP8;
    input wire n11XP2;
    input wire n1XP10;
    input wire n2XP3;
    input wire n2XP5;
    input wire n2XP7;
    input wire n2XP8;
    input wire n3XP2;
    input wire n3XP6;
    input wire n3XP7;
    input wire n4XP11;
    input wire n5XP12;
    input wire n5XP15;
    input wire n5XP21;
    input wire n5XP28;
    input wire n5XP4;
    input wire n6XP5;
    input wire n6XP8;
    output wire n7XP14;
    input wire n7XP19;
    input wire n7XP4;
    input wire n7XP9;
    inout wire n8PP4;
    input wire n8XP6;
    input wire n9XP1;
    input wire n9XP5;

    pullup R6001(NET_278);
    pullup R6002(A2X_n);
    pullup R6003(RB_n);
    pullup R6004(WYD_n);
    pullup R6005(NET_264);
    pullup R6006(WL_n);
    pullup R6007(RG_n);
    pullup R6008(WB_n);
    pullup R6009(RU_n);
    pullup R6010(WZ_n);
    pullup R6011(TOV_n);
    pullup R6012(WSC_n);
    pullup R6013(WG_n);
    pullup R6014(NET_255);
    pullup R6015(NET_219);
    pullup R6016(MONEX_n);
    pullup R6017(__A06_2__RB1_n);
    pullup R6018(__A06_2__R1C_n);
    pullup R6019(n8PP4);
    pullup R6020(NET_199);
    pullup R6021(WS_n);
    pullup R6022(NET_204);
    pullup R6023(CI_n);
    pullup R6024(WA_n);
    pullup R6025(NET_236);
    pullup R6026(ST2_n);
    pullup R6027(RZ_n);
    pullup R6028(RC_n);
    U74HC27 U6001(T04, T07, NET_281, NET_282, NET_283, NET_297, GND, NET_296, T01, T03, T05, NET_280, T10, VCC, SIM_RST);
    U74HC02 U6002(NET_281, NET_280, DV376_n, NET_282, T01_n, DV1376_n, GND, T04_n, DV4_n, NET_283, MP1_n, NET_278, NET_279, VCC, SIM_RST);
    U74HC27 U6003(T07, T09, L15A_n, L02A_n, L01_n, NET_295, GND, NET_311, T05, T08, T11, NET_294, T11, VCC, SIM_RST);
    U74LVC07 U6004(NET_296, NET_278, NET_294, NET_278, NET_305, A2X_n, GND, RB_n, NET_304, WYD_n, NET_306, WY_n, NET_301, VCC, SIM_RST);
    U74HC02 U6005(NET_330, NET_279, n2XP7, L2GD_n, __A06_1__ZIP, CGMC, GND, CGMC, NET_299, NET_306, NET_302, NET_298, NET_300, VCC, SIM_RST);
    U74HC04 U6006(L01_n, NET_293, L02A_n, NET_326, L15A_n, NET_331, GND, CGMC, NET_297, __A06_1__ZIP, NET_330, NET_328, NET_327, VCC, SIM_RST);
    U74HC27 U6007(n7XP19, __A06_1__ZIP, CGMC, NET_269, RBSQ, NET_304, GND, NET_307, NET_293, NET_326, NET_331, NET_305, CGMC, VCC, SIM_RST);
    U74HC27 U6008(NET_331, NET_293, NET_330, NET_298, NET_302, NET_301, GND, NET_327, NET_302, NET_298, L02A_n, NET_298, L02A_n, VCC, SIM_RST);
    U74HC02 U6009(NET_299, NET_330, NET_300, NET_303, NET_330, NET_328, GND, NET_311, DV376_n, NET_268, DV1376_n, T02_n, NET_329, VCC, SIM_RST);
    U74HC04 U6010(NET_303, __A06_1__MCRO_n, NET_273, NET_288, NET_271, NET_292, GND, __A06_1__ZAP, ZAP_n, NET_313, NET_311, __A06_1__MONEX, MONEX_n, VCC, SIM_RST);
    U74HC27 U6011(NET_330, NET_328, NET_327, NET_307, NET_330, NET_269, GND, NET_302, NET_326, L15A_n, L01_n, __A06_1__ZIPCI, NET_295, VCC, SIM_RST);
    U74HC02 U6012(NET_273, NET_268, NET_329, NET_271, NET_270, DIVSTG, GND, T08, T10, NET_262, MP1_n, NET_264, NET_267, VCC, SIM_RST);
    U74HC27 U6013(T06, T09, DV376_n, NET_272, T12USE_n, NET_270, GND, NET_263, T02, T04, T06, NET_272, T12, VCC, SIM_RST);
    U74LVC07 U6014(NET_263, NET_264, NET_262, NET_264, NET_287, WL_n, GND, RG_n, NET_284, WB_n, NET_289, RU_n, NET_277, VCC, SIM_RST);
    U74HC02 U6015(NET_266, T01, T03, NET_265, NET_266, MP3_n, GND, NET_267, NET_265, ZAP_n, n5XP28, NET_288, TSGU_n, VCC, SIM_RST);
    U74HC02 U6016(NET_287, NET_288, n5XP12, NET_274, RRPA, n5XP4, GND, n5XP15, n3XP6, WQ_n, n9XP5, n6XP8, NET_333, VCC, SIM_RST);
    U74HC4002 U6017(NET_284, n5XP4, RADRG, NET_288, n5XP28, NET_285, GND, NET_286, n5XP28, n1XP10, NET_292, n2XP3, NET_289, VCC, SIM_RST);
    U74HC4002 U6018(NET_277, NET_292, __A06_1__ZAP, n5XP12, n6XP5, NET_275, GND, NET_276, PRINC, DINC_n, MINC, DINC, NET_227, VCC, SIM_RST);
    U74LVC07 U6019(NET_274, WZ_n, NET_332, TOV_n, NET_333, WSC_n, GND, WG_n, NET_312, NET_255, NET_260, NET_255, NET_259, VCC, SIM_RST);
    U74HC27 U6020(n6XP5, n3XP2, BR1_n, PHS4_n, TSGU_n, __A06_1__RB1F, GND, __A06_1__CLXC, TSGU_n, BR1, PHS4_n, NET_332, n9XP5, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U6021(NET_312, n6XP8, n6XP8, PIFL_n, CGMC, NET_308, GND, PTWOX, __A06_1__MONEX, NET_310, __A06_1__MONEX, B15X, NET_309, VCC, SIM_RST);
    U74HC27 U6022(PIFL_n, NET_313, STBE, n1XP10, STBF, NET_315, GND, NET_260, NET_257, NET_256, INCR0, NET_308, T02, VCC, SIM_RST);
    U74HC04 U6023(NET_310, __A06_1__TWOX, NET_309, __A06_1__BXVX, NET_323, NET_324, GND, NET_325, NET_324, NET_322, NET_325, NET_319, NET_322, VCC, SIM_RST);
    U74HC02 U6024(__A06_1__CGMC, NET_315, NET_323, NET_321, __A06_1__CGMC, NET_314, GND, NET_321, NET_315, NET_323, BR1, AUG0_n, NET_257, VCC, SIM_RST);
    U74HC04 U6025(NET_319, NET_318, NET_318, NET_316, NET_316, NET_317, GND, NET_314, NET_317, NET_220, NET_218, NET_229, __A06_2__7XP10, VCC, SIM_RST);
    U74HC02 U6026(NET_256, DIM0_n, BR12B_n, NET_259, PINC, NET_258, GND, BR12B_n, DINC_n, NET_258, T06_n, NET_255, __A06_2__6XP10, VCC, SIM_RST);
    U74HC02 U6027(NET_214, MINC, MCDU, NET_212, AUG0_n, BR1_n, GND, DIM0_n, BR1B2B_n, NET_211, BR1B2B_n, DINC_n, NET_213, VCC, SIM_RST);
    U74HC27 U6028(NET_212, NET_211, BR1B2B_n, CDUSTB_n, DINC_n, __A06_2__POUT, GND, __A06_2__MOUT, BR12B_n, CDUSTB_n, DINC_n, NET_215, NET_213, VCC, SIM_RST);
    U74LVC07 U6029(NET_214, NET_219, NET_215, NET_219, NET_220, MONEX_n, GND, WA_n, NET_209, __A06_2__RB1_n, NET_229, __A06_2__R1C_n, NET_232, VCC, SIM_RST);
    U74HC02 U6030(NET_218, T06_n, NET_219, NET_216, PCDU, MCDU, GND, T06_n, NET_216, __A06_2__6XP12, NET_205, T07_n, NET_208, VCC, SIM_RST);
    U74HC27 U6031(BR2_n, DINC_n, DAS0, DAS1, MSU0, NET_205, GND, NET_209, NET_208, __A06_2__7XP7, NET_203, __A06_2__ZOUT, CDUSTB_n, VCC, SIM_RST);
    U74HC02 U6032(NET_210, DV4_n, BR1B2B, __A06_2__7XP7, T07_n, NET_206, GND, WAND0, INOTLD, NET_231, T07_n, NET_231, n7XP14, VCC, SIM_RST);
    U74HC27 U6033(NET_210, WAND0, DAS1_n, T07_n, BR1B2_n, __A06_2__7XP10, GND, __A06_2__7XP11, DAS1_n, T07_n, BR12B_n, NET_206, RAND0, VCC, SIM_RST);
    U74HC04 U6034(__A06_2__7XP11, NET_232, NET_190, __A06_2__PONEX, ST2_n, ST2, GND, ST1, NET_245, NET_242, __A06_2__PSEUDO, NET_243, __A06_2__RDBANK, VCC, SIM_RST);
    U74HC02 U6035(__A06_2__7XP15, NET_223, T07_n, NET_226, NET_227, T07_n, GND, PRINC, INKL, NET_225, IC9, DXCH0, NET_187, VCC, SIM_RST);
    U74HC27 U6036(PCDU, MCDU, n7XP9, n11XP2, __A06_2__7XP15, RUS_n, GND, NET_228, NET_226, NET_234, NET_203, NET_223, SHIFT, VCC, SIM_RST);
    U74LVC07 U6037(NET_228, RU_n, NET_183, WSC_n, NET_184, WG_n, GND, RB_n, NET_186, n8PP4, NET_179, n8PP4, NET_177, VCC, SIM_RST);
    U74HC27 U6038(NET_225, T07_n, T04_n, MON_n, FETCH1, NET_185, GND, NET_183, __A06_2__WOVR, NET_185, NET_240, __A06_2__WOVR, MONPCH, VCC, SIM_RST);
    U74HC02 U6039(NET_184, __A06_2__WOVR, NET_240, NET_240, T07_n, NET_187, GND, __A06_2__10XP9, NET_240, NET_186, T08_n, n8PP4, __A06_2__8XP4, VCC, SIM_RST);
    U74HC27 U6040(RUPT1, DAS1, IC17, MASK0, IC11, NET_177, GND, NET_178, IC6, IC7, DV4B1B, NET_179, DV4_n, VCC, SIM_RST);
    U74LVC07 U6041(NET_178, n8PP4, NET_181, NET_199, NET_180, NET_199, GND, WS_n, NET_200, NET_204, NET_198, NET_204, NET_201, VCC, SIM_RST);
    U74HC27 U6042(T08_n, RUPT0, NET_199, R6, R15, NET_200, GND, NET_201, ADS0, IC11, NET_202, NET_181, DAS0, VCC, SIM_RST);
    U74HC02 U6043(NET_180, MP1, DV1376, NET_197, MP3_n, BR1_n, GND, NET_197, CCS0, NET_198, T11_n, NET_204, NET_203, VCC, SIM_RST);
    U74HC02 U6044(NET_202, DAS1_n, BR2_n, NET_189, __A06_1__ZIPCI, __A06_2__6XP12, GND, CCS0_n, BR1B2B_n, NET_195, T10_n, NDXX1_n, EXT, VCC, SIM_RST);
    U74HC27 U6045(T03_n, DAS1_n, NET_239, NET_234, n2XP5, NET_253, GND, NET_248, IC7, DCS0, SU0, NET_234, ADS0, VCC, SIM_RST);
    U74HC4002 U6046(NET_190, n8XP6, n7XP4, n10XP8, __A06_2__6XP10, NET_191, GND, NET_192, IC6, DCA0, AD0, NET_195, NET_196, VCC, SIM_RST);
    U74LVC07 U6047(NET_189, CI_n, NET_253, WA_n, NET_254, RC_n, GND, NET_236, NET_248, NET_236, NET_249, ST2_n, NET_252, VCC, SIM_RST);
    U74HC02 U6048(__A06_2__10XP9, T10_n, NET_196, NET_238, IC6, IC7, GND, T10_n, NET_238, NET_239, T10_n, NET_236, NET_235, VCC, SIM_RST);
    U74HC02 U6049(NET_254, NET_235, __A06_2__7XP7, NET_249, NET_237, DV4B1B, GND, CCS0_n, BR12B_n, NET_237, T10_n, MP1_n, __A06_2__10XP15, VCC, SIM_RST);
    U74HC27 U6050(__A06_2__8XP4, __A06_2__10XP15, __A06_2__8XP4, RADRZ, n9XP1, NET_244, GND, NEAC, NET_246, TL15, GOJAM, NET_252, RADRZ, VCC, SIM_RST);
    wire U6051_9_NC;
    wire U6051_10_NC;
    wire U6051_11_NC;
    wire U6051_12_NC;
    wire U6051_13_NC;
    U74HC4002 U6051(NET_245, n2XP8, n10XP1, MP0T10, __A06_2__10XP15, NET_250, GND, NET_251, U6051_9_NC, U6051_10_NC, U6051_11_NC, U6051_12_NC, U6051_13_NC, VCC, SIM_RST);
    wire U6052_10_NC;
    wire U6052_11_NC;
    wire U6052_12_NC;
    wire U6052_13_NC;
    U74LVC07 U6052(NET_244, RZ_n, NET_242, RPTSET, NET_243, RU_n, GND, RC_n, NET_320, U6052_10_NC, U6052_11_NC, U6052_12_NC, U6052_13_NC, VCC, SIM_RST);
    U74HC02 #(1, 0, 0, 0) U6053(NET_246, MP0T10, NEAC, NET_241, RADRZ, __A06_2__PSEUDO, GND, T06_n, STFET1_n, __A06_2__RDBANK, __A06_1__ZIPCI, n3XP7, NET_320, VCC, SIM_RST);
    wire U6054_8_NC;
    wire U6054_9_NC;
    wire U6054_10_NC;
    wire U6054_11_NC;
    U74HC27 #(1, 0, 0) U6054(NET_241, GOJAM, n3XP7, n5XP21, n4XP11, RCH_n, GND, U6054_8_NC, U6054_9_NC, U6054_10_NC, U6054_11_NC, __A06_2__PSEUDO, RADRG, VCC, SIM_RST);
endmodule