`include "components/agc_parts.v"

module stage_branch(VCC, GND, SIM_RST, GOJAM, T01, T03, T12_n, PHS3_n, ST1, ST2, INKL, STRTFC, DVST, DVST_n, RSTSTG, TRSM_n, XT1_n, XB7_n, NDR100_n, ST0_n, ST1_n, STD2, ST3_n, ST4, MTCSAI);
    input wire SIM_RST;
    input wire DVST;
    input wire DVST_n;
    input wire GND;
    input wire GOJAM;
    input wire INKL;
    input wire MTCSAI;
    input wire NDR100_n;
    wire NET_34;
    wire NET_35;
    wire NET_36;
    wire NET_37;
    wire NET_38;
    wire NET_41;
    wire NET_42;
    wire NET_43;
    wire NET_44;
    wire NET_45;
    wire NET_46;
    wire NET_47;
    wire NET_48;
    wire NET_49;
    wire NET_50;
    wire NET_51;
    wire NET_52;
    wire NET_53;
    wire NET_54;
    wire NET_55;
    wire NET_56;
    wire NET_57;
    wire NET_58;
    wire NET_59;
    wire NET_60;
    wire NET_61;
    wire NET_62;
    wire NET_63;
    wire NET_64;
    wire NET_65;
    wire NET_66;
    wire NET_67;
    wire NET_68;
    wire NET_69;
    wire NET_70;
    input wire PHS3_n;
    input wire RSTSTG;
    output wire ST0_n;
    input wire ST1;
    output wire ST1_n;
    input wire ST2;
    output wire ST3_n;
    input wire ST4;
    wire ST4_n;
    output wire STD2;
    input wire STRTFC;
    input wire T01;
    input wire T03;
    input wire T12_n;
    input wire TRSM_n;
    input wire VCC;
    input wire XB7_n;
    input wire XT1_n;
    wire __A04_1__DIVSTG;
    wire __A04_1__MST1;
    wire __A04_1__MST2;
    wire __A04_1__MST3;
    wire __A04_1__STG1;
    wire __A04_1__STG2;
    wire __A04_1__STG3;
    wire __A04_1__T12USE_n;

    pullup R4001(NET_55);
    pullup R4002(NET_62);
    U74HC02 #(0, 0, 0, 1) U4001(__A04_1__T12USE_n, DVST, NET_59, __A04_1__DIVSTG, __A04_1__T12USE_n, T03, GND, NET_58, NET_60, NET_70, GOJAM, MTCSAI, NET_54, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U4002(T03, __A04_1__T12USE_n, __A04_1__T12USE_n, RSTSTG, GOJAM, NET_59, GND, NET_60, PHS3_n, NET_59, T12_n, NET_58, PHS3_n, VCC, SIM_RST);
    wire U4003_10_NC;
    wire U4003_11_NC;
    wire U4003_12_NC;
    wire U4003_13_NC;
    U74LVC07 U4003(NET_54, NET_55, NET_57, NET_55, NET_61, NET_62, GND, NET_62, NET_67, U4003_10_NC, U4003_11_NC, U4003_12_NC, U4003_13_NC, VCC, SIM_RST);
    U74HC27 #(1, 1, 0) U4004(ST1, NET_56, __A04_1__STG1, __A04_1__STG3, __A04_1__STG2, NET_65, GND, NET_64, __A04_1__STG2, __A04_1__STG3, NET_34, NET_57, NET_44, VCC, SIM_RST);
    U74HC02 U4005(NET_44, NET_55, T01, NET_56, DVST_n, NET_52, GND, NET_70, NET_55, NET_69, NET_44, NET_70, NET_68, VCC, SIM_RST);
    U74HC02 #(1, 0, 1, 0) U4006(NET_34, NET_69, __A04_1__STG1, __A04_1__STG1, NET_34, NET_68, GND, ST2, NET_42, NET_61, DVST_n, NET_34, NET_63, VCC, SIM_RST);
    wire U4007_8_NC;
    wire U4007_9_NC;
    wire U4007_10_NC;
    wire U4007_11_NC;
    wire U4007_12_NC;
    wire U4007_13_NC;
    U74HC04 U4007(NET_34, __A04_1__MST1, NET_38, __A04_1__MST2, NET_52, __A04_1__MST3, GND, U4007_8_NC, U4007_9_NC, U4007_10_NC, U4007_11_NC, U4007_12_NC, U4007_13_NC, VCC, SIM_RST);
    wire U4008_10_NC;
    wire U4008_11_NC;
    wire U4008_12_NC;
    wire U4008_13_NC;
    U74HC04 #(0, 1, 1, 1, 0, 0) U4008(NET_65, ST0_n, NET_64, ST1_n, NET_45, ST3_n, GND, ST4_n, NET_48, U4008_10_NC, U4008_11_NC, U4008_12_NC, U4008_13_NC, VCC, SIM_RST);
    U74HC27 #(1, 0, 0) U4009(NET_63, MTCSAI, NET_62, GOJAM, T01, NET_66, GND, NET_45, __A04_1__STG3, NET_38, NET_34, NET_67, NET_66, VCC, SIM_RST);
    U74HC4002 U4010(NET_42, TRSM_n, XT1_n, XB7_n, NDR100_n, NET_41, GND, NET_43, NET_50, STRTFC, T01, RSTSTG, NET_49, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U4011(NET_36, NET_70, NET_62, NET_35, NET_66, NET_70, GND, NET_36, __A04_1__STG2, NET_38, NET_38, NET_35, __A04_1__STG2, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U4012(NET_37, DVST_n, NET_38, NET_50, NET_37, NET_49, GND, NET_70, NET_50, NET_51, NET_49, NET_70, NET_53, VCC, SIM_RST);
    wire U4013_8_NC;
    wire U4013_9_NC;
    wire U4013_10_NC;
    wire U4013_11_NC;
    wire U4013_12_NC;
    wire U4013_13_NC;
    U74HC02 #(1, 0, 0, 0) U4013(NET_52, NET_51, __A04_1__STG3, __A04_1__STG3, NET_52, NET_53, GND, U4013_8_NC, U4013_9_NC, U4013_10_NC, U4013_11_NC, U4013_12_NC, U4013_13_NC, VCC, SIM_RST);
    wire U4014_9_NC;
    wire U4014_10_NC;
    wire U4014_11_NC;
    wire U4014_12_NC;
    wire U4014_13_NC;
    U74HC4002 U4014(STD2, INKL, __A04_1__STG1, __A04_1__STG3, NET_38, NET_46, GND, NET_47, U4014_9_NC, U4014_10_NC, U4014_11_NC, U4014_12_NC, U4014_13_NC, VCC, SIM_RST);
    wire U4015_3_NC;
    wire U4015_4_NC;
    wire U4015_5_NC;
    wire U4015_6_NC;
    wire U4015_8_NC;
    wire U4015_9_NC;
    wire U4015_10_NC;
    wire U4015_11_NC;
    U74HC27 U4015(NET_52, __A04_1__STG1, U4015_3_NC, U4015_4_NC, U4015_5_NC, U4015_6_NC, GND, U4015_8_NC, U4015_9_NC, U4015_10_NC, U4015_11_NC, NET_48, __A04_1__STG2, VCC, SIM_RST);
endmodule