`timescale 1ns/1ps
`default_nettype none

module inout_vi(VCC, GND, SIM_RST, SIM_CLK, P04_n, SB2_n, F18A, F18B, F5ASB0_n, F5ASB2, F5ASB2_n, CCHG_n, WCHG_n, CCH11, CCH12, CCH13, CCH14, CCH33, RCH11_n, RCH12_n, RCH13_n, RCH14_n, WCH11_n, WCH12_n, WCH13_n, WCH14_n, POUT_n, MOUT_n, ZOUT_n, T6RPT, PIPPLS_n, PIPAXp, PIPAXm, PIPAYp, PIPAYm, PIPAZp, PIPAZm, OCTAD5, CHWL05_n, CHWL06_n, CHWL07_n, CHWL08_n, CHWL10_n, CHWL11_n, CHWL12_n, CHWL13_n, CHWL14_n, CHWL16_n, XT0_n, XB0_n, XB1_n, XB2_n, XB3_n, XB4_n, XB7_n, T6ON_n, ALTEST, E5, E6, E7_n, CDUXD, CDUYD, CDUZD, PIPAFL, PIPXP, PIPXM, PIPYP, PIPYM, PIPZP, PIPZM, TRUND, SHAFTD, CH0705, CH0706, CH0707, CH1310, CH1316, CH1411, CH1412, CH1413, CH1414, CH1416, CH1108, CH1113, CH1114, CH1116, CH1216, CDUXDP, CDUXDM, CDUYDP, CDUYDM, CDUZDP, CDUZDM);
    input wire VCC;
    input wire GND;
    input wire SIM_RST;
    input wire SIM_CLK;
    output wire ALTEST;
    input wire CCH11;
    input wire CCH12;
    input wire CCH13;
    input wire CCH14;
    input wire CCH33;
    input wire CCHG_n;
    output wire CDUXD;
    output wire CDUXDM;
    output wire CDUXDP;
    output wire CDUYD;
    output wire CDUYDM;
    output wire CDUYDP;
    output wire CDUZD;
    output wire CDUZDM;
    output wire CDUZDP;
    output wire CH0705;
    output wire CH0706;
    output wire CH0707;
    output wire CH1108;
    output wire CH1113;
    output wire CH1114;
    output wire CH1116;
    output wire CH1216;
    output wire CH1310;
    output wire CH1316;
    output wire CH1411;
    output wire CH1412;
    output wire CH1413;
    output wire CH1414;
    output wire CH1416;
    input wire CHWL05_n;
    input wire CHWL06_n;
    input wire CHWL07_n;
    input wire CHWL08_n;
    input wire CHWL10_n;
    input wire CHWL11_n;
    input wire CHWL12_n;
    input wire CHWL13_n;
    input wire CHWL14_n;
    input wire CHWL16_n;
    output wire E5;
    output wire E6;
    output wire E7_n;
    input wire F18A;
    input wire F18B;
    input wire F5ASB0_n;
    input wire F5ASB2;
    input wire F5ASB2_n;
    input wire MOUT_n;
    input wire OCTAD5;
    input wire P04_n;
    output wire PIPAFL;
    input wire PIPAXm;
    input wire PIPAXp;
    input wire PIPAYm;
    input wire PIPAYp;
    input wire PIPAZm;
    input wire PIPAZp;
    input wire PIPPLS_n;
    output wire PIPXM;
    output wire PIPXP;
    output wire PIPYM;
    output wire PIPYP;
    output wire PIPZM;
    output wire PIPZP;
    input wire POUT_n;
    input wire RCH11_n;
    input wire RCH12_n;
    input wire RCH13_n;
    input wire RCH14_n;
    input wire SB2_n;
    output wire SHAFTD;
    output wire T6ON_n;
    input wire T6RPT;
    output wire TRUND;
    input wire WCH11_n;
    input wire WCH12_n;
    input wire WCH13_n;
    input wire WCH14_n;
    input wire WCHG_n;
    input wire XB0_n;
    input wire XB1_n;
    input wire XB2_n;
    input wire XB3_n;
    input wire XB4_n;
    input wire XB7_n;
    input wire XT0_n;
    input wire ZOUT_n;
    wire __A23_1__BOTHX;
    wire __A23_1__BOTHY;
    wire __A23_1__BOTHZ;
    wire __A23_1__F18AX;
    wire __A23_1__F18A_n;
    wire __A23_1__F18B_n;
    wire __A23_1__MISSX;
    wire __A23_1__MISSY;
    wire __A23_1__MISSZ;
    wire __A23_1__NOXM;
    wire __A23_1__NOXP;
    wire __A23_1__NOYM;
    wire __A23_1__NOYP;
    wire __A23_1__NOZM;
    wire __A23_1__NOZP;
    wire __A23_1__P04A;
    wire __A23_1__PIPAXm_n;
    wire __A23_1__PIPAXp_n;
    wire __A23_1__PIPAYm_n;
    wire __A23_1__PIPAYp_n;
    wire __A23_1__PIPAZm_n;
    wire __A23_1__PIPAZp_n;
    wire __A23_1__PIPGXm;
    wire __A23_1__PIPGXp;
    wire __A23_1__PIPGYm;
    wire __A23_1__PIPGYp;
    wire __A23_1__PIPGZm;
    wire __A23_1__PIPGZp;
    wire __A23_1__PIPSAM;
    wire __A23_1__PIPSAM_n;
    wire __A23_2__CCH07;
    wire __A23_2__ISSTDC;
    wire __A23_2__OT1108;
    wire __A23_2__OT1113;
    wire __A23_2__OT1114;
    wire __A23_2__OT1116;
    wire __A23_2__RCH07_n;
    wire __A23_2__SHFTDM;
    wire __A23_2__SHFTDP;
    wire __A23_2__TRNDM;
    wire __A23_2__TRNDP;
    wire __A23_2__WCH07_n;
    wire __A23_NET_101;
    wire __A23_NET_102;
    wire __A23_NET_103;
    wire __A23_NET_104;
    wire __A23_NET_105;
    wire __A23_NET_106;
    wire __A23_NET_107;
    wire __A23_NET_108;
    wire __A23_NET_109;
    wire __A23_NET_110;
    wire __A23_NET_111;
    wire __A23_NET_112;
    wire __A23_NET_113;
    wire __A23_NET_114;
    wire __A23_NET_115;
    wire __A23_NET_116;
    wire __A23_NET_117;
    wire __A23_NET_118;
    wire __A23_NET_120;
    wire __A23_NET_121;
    wire __A23_NET_124;
    wire __A23_NET_125;
    wire __A23_NET_126;
    wire __A23_NET_127;
    wire __A23_NET_128;
    wire __A23_NET_129;
    wire __A23_NET_130;
    wire __A23_NET_132;
    wire __A23_NET_147;
    wire __A23_NET_149;
    wire __A23_NET_151;
    wire __A23_NET_153;
    wire __A23_NET_154;
    wire __A23_NET_157;
    wire __A23_NET_158;
    wire __A23_NET_159;
    wire __A23_NET_160;
    wire __A23_NET_161;
    wire __A23_NET_162;
    wire __A23_NET_164;
    wire __A23_NET_165;
    wire __A23_NET_166;
    wire __A23_NET_168; //FPGA#wand
    wire __A23_NET_170;
    wire __A23_NET_171;
    wire __A23_NET_172;
    wire __A23_NET_173;
    wire __A23_NET_174;
    wire __A23_NET_175;
    wire __A23_NET_176;
    wire __A23_NET_177;
    wire __A23_NET_178;
    wire __A23_NET_179;
    wire __A23_NET_180;
    wire __A23_NET_181;
    wire __A23_NET_182;
    wire __A23_NET_185;
    wire __A23_NET_186;
    wire __A23_NET_187;
    wire __A23_NET_188;
    wire __A23_NET_189; //FPGA#wand
    wire __A23_NET_190;
    wire __A23_NET_191;
    wire __A23_NET_192;
    wire __A23_NET_193;
    wire __A23_NET_194;
    wire __A23_NET_195;
    wire __A23_NET_196;
    wire __A23_NET_197;
    wire __A23_NET_198;
    wire __A23_NET_199;
    wire __A23_NET_200;
    wire __A23_NET_201;
    wire __A23_NET_202;
    wire __A23_NET_203;
    wire __A23_NET_205;
    wire __A23_NET_206;
    wire __A23_NET_207;
    wire __A23_NET_208;
    wire __A23_NET_209;
    wire __A23_NET_210;
    wire __A23_NET_212;
    wire __A23_NET_213;
    wire __A23_NET_214;
    wire __A23_NET_215;
    wire __A23_NET_216;
    wire __A23_NET_217;
    wire __A23_NET_218;
    wire __A23_NET_219;
    wire __A23_NET_220;
    wire __A23_NET_221;
    wire __A23_NET_222;
    wire __A23_NET_223;
    wire __A23_NET_227;
    wire __A23_NET_228;
    wire __A23_NET_229;
    wire __A23_NET_230;
    wire __A23_NET_231;
    wire __A23_NET_232;
    wire __A23_NET_233;
    wire __A23_NET_234;
    wire __A23_NET_235;
    wire __A23_NET_236;
    wire __A23_NET_237;
    wire __A23_NET_238;
    wire __A23_NET_239;
    wire __A23_NET_240;
    wire __A23_NET_241;
    wire __A23_NET_242;
    wire __A23_NET_243;
    wire __A23_NET_244;
    wire __A23_NET_245;
    wire __A23_NET_246;
    wire __A23_NET_247;
    wire __A23_NET_248;
    wire __A23_NET_249;
    wire __A23_NET_250;
    wire __A23_NET_251;
    wire __A23_NET_252;
    wire __A23_NET_253;
    wire __A23_NET_254;
    wire __A23_NET_255;
    wire __A23_NET_256;
    wire __A23_NET_257;
    wire __A23_NET_258;
    wire __A23_NET_259;
    wire __A23_NET_260;
    wire __A23_NET_261;
    wire __A23_NET_262;
    wire __A23_NET_263;
    wire __A23_NET_264;
    wire __A23_NET_265;
    wire __A23_NET_266;
    wire __A23_NET_267;
    wire __A23_NET_268;
    wire __A23_NET_269;
    wire __A23_NET_270;
    wire __A23_NET_271;
    wire __A23_NET_272;
    wire __A23_NET_273;

    pullup R23001(__A23_NET_168);
    pullup R23002(__A23_NET_189);
    U74HC27 #(1'b1, 1'b1, 1'b1) U23001(__A23_1__NOXP, __A23_1__NOXM, __A23_1__NOYM, __A23_1__NOZP, __A23_1__NOZM, __A23_NET_188, GND, __A23_NET_166, __A23_1__MISSX, __A23_1__MISSY, __A23_1__MISSZ, __A23_NET_187, __A23_1__NOYP, VCC, SIM_RST, SIM_CLK);
    U74LVC07 U23002(__A23_NET_187, __A23_NET_168, __A23_NET_188, __A23_NET_168, __A23_NET_185, __A23_NET_189, GND, __A23_NET_189, __A23_NET_186,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK); //FPGA#OD:2,4,6,8
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1) U23003(F18B, __A23_1__F18B_n, __A23_1__PIPGXp, __A23_NET_209, __A23_1__PIPGXm, __A23_NET_208, GND, __A23_NET_160, F5ASB2, __A23_NET_129, __A23_1__PIPGYp, __A23_NET_130, __A23_1__PIPGYm, VCC, SIM_RST, SIM_CLK);
    U74HC02 U23004(__A23_NET_164, __A23_1__F18B_n, __A23_NET_168, __A23_NET_165, F5ASB0_n, __A23_NET_166, GND, __A23_NET_189, CCH33, PIPAFL, __A23_NET_172, __A23_NET_170, __A23_NET_161, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b1, 1'b0) U23005(__A23_1__BOTHX, __A23_1__BOTHY, __A23_NET_164, __A23_NET_165, PIPAFL, __A23_NET_186, GND, __A23_NET_171, __A23_NET_173, __A23_NET_207, __A23_NET_209, __A23_NET_185, __A23_1__BOTHZ, VCC, SIM_RST, SIM_CLK);
    U74HC27 U23006(__A23_NET_208, __A23_NET_207,  ,  ,  ,  , GND,  ,  ,  ,  , __A23_NET_172, __A23_NET_162, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23007(__A23_NET_170, __A23_NET_161, __A23_NET_171, __A23_NET_158, __A23_NET_160, __A23_NET_161, GND, __A23_NET_170, __A23_NET_160, __A23_NET_159, __A23_NET_158, __A23_NET_162, __A23_NET_173, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23008(__A23_NET_162, __A23_NET_173, __A23_NET_159, __A23_NET_182, __A23_NET_160, __A23_NET_179, GND, __A23_NET_174, __A23_NET_160, __A23_NET_180, __A23_NET_182, __A23_NET_207, __A23_NET_181, VCC, SIM_RST, SIM_CLK);
    U74HC27 U23009(__A23_NET_162, __A23_NET_207, __A23_NET_173, __A23_NET_207, __A23_NET_208, __A23_NET_175, GND, __A23_NET_178, __A23_NET_162, __A23_NET_181, __A23_NET_208, __A23_NET_176, __A23_NET_209, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U23010(__A23_NET_173, __A23_NET_181, __A23_NET_176, __A23_NET_175, __A23_NET_174, __A23_NET_179, GND, __A23_NET_174, __A23_NET_179, __A23_NET_178, __A23_NET_177, __A23_NET_177, __A23_NET_209, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U23011(__A23_NET_207, __A23_NET_181, __A23_NET_180, __A23_1__BOTHX, __A23_NET_208, __A23_NET_209, GND, __A23_1__PIPGXm, __A23_NET_205, __A23_1__NOXM, __A23_1__NOXM, __A23_1__F18AX, __A23_NET_205, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23012(__A23_1__NOXP, __A23_1__PIPGXp, __A23_NET_206, __A23_NET_206, __A23_1__NOXP, __A23_1__F18AX, GND, __A23_1__MISSX, F5ASB2, __A23_NET_210, __A23_NET_130, __A23_NET_129, __A23_1__BOTHY, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U23013(__A23_1__PIPGXp, __A23_1__PIPGXm, __A23_NET_162, __A23_NET_181, __A23_NET_209, PIPXP, GND, PIPXM, __A23_NET_173, __A23_NET_181, __A23_NET_208, __A23_1__MISSX, __A23_NET_210, VCC, SIM_RST, SIM_CLK);
    U74HC27 U23014(__A23_NET_130, __A23_NET_202, __A23_NET_128, __A23_NET_202, __A23_NET_129, __A23_NET_190, GND, __A23_NET_126, __A23_NET_196, __A23_NET_202, __A23_NET_129, __A23_NET_193, __A23_NET_196, VCC, SIM_RST, SIM_CLK);
    U74HC27 U23015(__A23_NET_128, __A23_NET_202, __A23_NET_196, __A23_NET_201, __A23_NET_130, __A23_NET_125, GND, __A23_NET_124, __A23_NET_128, __A23_NET_201, __A23_NET_129, __A23_NET_127, __A23_NET_130, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23016(__A23_NET_191, __A23_NET_193, __A23_NET_192, __A23_NET_192, __A23_NET_191, __A23_NET_190, GND, __A23_NET_203, __A23_NET_191, __A23_NET_195, __A23_NET_192, __A23_NET_203, __A23_NET_194, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b1) U23017(__A23_NET_126, __A23_NET_127, __A23_NET_197, __A23_NET_125, __A23_NET_124, __A23_NET_198, GND, __A23_1__MISSY, __A23_1__PIPGYp, __A23_1__PIPGYm, __A23_NET_132, __A23_NET_197, __A23_NET_198, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0) U23018(F5ASB2, __A23_NET_203, __A23_1__PIPGZp, __A23_NET_147, __A23_1__PIPGZm, __A23_NET_104, GND, __A23_NET_102, F5ASB2, __A23_1__F18A_n, F18A, __A23_1__F18AX, __A23_1__F18A_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U23019(__A23_NET_199, __A23_NET_203, __A23_NET_197, __A23_NET_200, __A23_NET_198, __A23_NET_203, GND, __A23_NET_195, __A23_NET_196, __A23_NET_128, __A23_NET_128, __A23_NET_194, __A23_NET_196, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U23020(__A23_NET_201, __A23_NET_199, __A23_NET_202, __A23_NET_202, __A23_NET_201, __A23_NET_200, GND, __A23_1__PIPGYm, __A23_NET_120, __A23_1__NOYM, __A23_1__NOYM, __A23_1__F18AX, __A23_NET_120, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23021(__A23_1__NOYP, __A23_1__PIPGYp, __A23_NET_121, __A23_NET_121, __A23_1__NOYP, __A23_1__F18AX, GND, __A23_1__MISSY, F5ASB2, __A23_NET_132, __A23_NET_104, __A23_NET_147, __A23_1__BOTHZ, VCC, SIM_RST, SIM_CLK);
    U74HC27 U23022(__A23_NET_196, __A23_NET_201, __A23_NET_128, __A23_NET_201, __A23_NET_130, PIPYM, GND, __A23_NET_107, __A23_NET_104, __A23_NET_151, __A23_NET_101, PIPYP, __A23_NET_129, VCC, SIM_RST, SIM_CLK);
    U74HC27 U23023(__A23_NET_108, __A23_NET_151, __A23_NET_101, __A23_NET_151, __A23_NET_147, __A23_NET_116, GND, __A23_NET_115, __A23_NET_108, __A23_NET_151, __A23_NET_104, __A23_NET_106, __A23_NET_147, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U23024(__A23_NET_101, __A23_NET_154, __A23_NET_108, __A23_NET_154, __A23_NET_147, __A23_NET_117, GND, __A23_1__MISSZ, __A23_1__PIPGZp, __A23_1__PIPGZm, __A23_NET_153, __A23_NET_118, __A23_NET_104, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U23025(__A23_NET_103, __A23_NET_107, __A23_NET_105, __A23_NET_105, __A23_NET_103, __A23_NET_106, GND, __A23_1__PIPGZm, __A23_NET_149, __A23_1__NOZM, __A23_1__NOZM, __A23_1__F18AX, __A23_NET_149, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U23026(__A23_NET_116, __A23_NET_115, __A23_NET_113, __A23_NET_118, __A23_NET_117, __A23_NET_114, GND, PIPZP, __A23_NET_101, __A23_NET_154, __A23_NET_147, __A23_NET_113, __A23_NET_114, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23027(__A23_1__NOZP, __A23_1__PIPGZp, __A23_NET_157, __A23_NET_157, __A23_1__NOZP, __A23_1__F18AX, GND, __A23_1__MISSZ, F5ASB2, __A23_NET_153, __A23_NET_102, __A23_NET_103, __A23_NET_109, VCC, SIM_RST, SIM_CLK);
    U74HC02 U23028(__A23_NET_110, __A23_NET_105, __A23_NET_102, __A23_NET_111, __A23_NET_102, __A23_NET_113, GND, __A23_NET_114, __A23_NET_102, __A23_NET_112, __A23_NET_109, __A23_NET_101, __A23_NET_108, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U23029(__A23_NET_101, __A23_NET_108, __A23_NET_110, __A23_NET_154, __A23_NET_111, __A23_NET_151, GND, __A23_NET_154, __A23_NET_112, __A23_NET_151, CHWL16_n, WCH14_n, __A23_NET_253, VCC, SIM_RST, SIM_CLK);
    U74HC27 U23030(__A23_NET_108, __A23_NET_154, __A23_NET_255, CCH14, __A23_NET_256, __A23_NET_254, GND, __A23_NET_251, __A23_NET_246, CCH14, __A23_NET_244, PIPZM, __A23_NET_104, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23031(__A23_NET_255, __A23_NET_253, __A23_NET_254, CH1416, RCH14_n, __A23_NET_255, GND, __A23_NET_255, F5ASB2_n, CDUXD, XB0_n, __A23_NET_270, __A23_NET_252, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0) U23032(__A23_NET_252, __A23_NET_258, OCTAD5, __A23_NET_270, __A23_NET_243, __A23_NET_245, GND, __A23_NET_268, __A23_NET_267, __A23_NET_271, __A23_NET_269, __A23_NET_263, __A23_NET_264, VCC, SIM_RST, SIM_CLK);
    U74HC02 U23034(CDUXDP, POUT_n, __A23_NET_258, CDUXDM, MOUT_n, __A23_NET_258, GND, ZOUT_n, __A23_NET_258, __A23_NET_256, CHWL14_n, WCH14_n, __A23_NET_257, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23035(__A23_NET_246, __A23_NET_257, __A23_NET_251, CH1414, RCH14_n, __A23_NET_246, GND, __A23_NET_246, F5ASB2_n, CDUYD, XB1_n, __A23_NET_270, __A23_NET_243, VCC, SIM_RST, SIM_CLK);
    U74HC02 U23036(CDUYDP, POUT_n, __A23_NET_245, CDUYDM, MOUT_n, __A23_NET_245, GND, ZOUT_n, __A23_NET_245, __A23_NET_244, CHWL13_n, WCH14_n, __A23_NET_249, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23037(__A23_NET_250, __A23_NET_249, __A23_NET_248, CH1413, RCH14_n, __A23_NET_250, GND, __A23_NET_250, F5ASB2_n, CDUZD, XB2_n, __A23_NET_270, __A23_NET_267, VCC, SIM_RST, SIM_CLK);
    U74HC27 U23038(__A23_NET_250, CCH14, __A23_NET_273, CCH14, __A23_NET_262, __A23_NET_272, GND, __A23_NET_260, __A23_NET_265, CCH14, __A23_NET_261, __A23_NET_248, __A23_NET_247, VCC, SIM_RST, SIM_CLK);
    U74HC02 U23039(CDUZDP, POUT_n, __A23_NET_268, CDUZDM, MOUT_n, __A23_NET_268, GND, ZOUT_n, __A23_NET_268, __A23_NET_247, CHWL12_n, WCH14_n, __A23_NET_266, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23040(__A23_NET_273, __A23_NET_266, __A23_NET_272, CH1412, RCH14_n, __A23_NET_273, GND, __A23_NET_273, F5ASB2_n, TRUND, XB3_n, __A23_NET_270, __A23_NET_269, VCC, SIM_RST, SIM_CLK);
    U74HC02 U23041(__A23_2__TRNDP, POUT_n, __A23_NET_271, __A23_2__TRNDM, MOUT_n, __A23_NET_271, GND, ZOUT_n, __A23_NET_271, __A23_NET_262, CHWL11_n, WCH14_n, __A23_NET_259, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23042(__A23_NET_265, __A23_NET_259, __A23_NET_260, CH1411, RCH14_n, __A23_NET_265, GND, __A23_NET_265, F5ASB2_n, SHAFTD, XB4_n, __A23_NET_270, __A23_NET_264, VCC, SIM_RST, SIM_CLK);
    U74HC02 U23043(__A23_2__SHFTDP, POUT_n, __A23_NET_263, __A23_2__SHFTDM, MOUT_n, __A23_NET_263, GND, ZOUT_n, __A23_NET_263, __A23_NET_261, CHWL05_n, __A23_2__WCH07_n, __A23_NET_221, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23044(__A23_NET_222, __A23_NET_221, E5, E5, __A23_NET_222, __A23_2__CCH07, GND, __A23_2__RCH07_n, __A23_NET_222, CH0705, CHWL06_n, __A23_2__WCH07_n, __A23_NET_219, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23045(__A23_NET_220, __A23_NET_219, E6, E6, __A23_NET_220, __A23_2__CCH07, GND, __A23_2__RCH07_n, __A23_NET_220, CH0706, CHWL07_n, __A23_2__WCH07_n, __A23_NET_227, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23046(E7_n, __A23_NET_227, __A23_NET_223, __A23_NET_223, E7_n, __A23_2__CCH07, GND, __A23_2__RCH07_n, E7_n, CH0707, XB7_n, XT0_n, __A23_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC27 U23047(WCHG_n, XT0_n, CCHG_n, XB7_n, XT0_n, __A23_2__CCH07, GND, __A23_NET_228, T6ON_n, T6RPT, CCH13, __A23_NET_215, XB7_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U23048(__A23_NET_215, __A23_2__WCH07_n, __A23_NET_212, __A23_2__RCH07_n, __A23_NET_218, __A23_2__OT1108, GND, __A23_2__OT1113, __A23_NET_239, __A23_2__OT1114, __A23_NET_238, __A23_2__OT1116, __A23_NET_242, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23049(__A23_NET_214, CHWL08_n, WCH11_n, __A23_NET_218, __A23_NET_214, __A23_NET_213, GND, __A23_NET_218, CCH11, __A23_NET_213, RCH11_n, __A23_NET_218, CH1108, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23050(__A23_NET_217, CHWL13_n, WCH11_n, __A23_NET_239, __A23_NET_217, __A23_NET_216, GND, __A23_NET_239, CCH11, __A23_NET_216, RCH11_n, __A23_NET_239, CH1113, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23051(__A23_NET_236, CHWL14_n, WCH11_n, __A23_NET_238, __A23_NET_236, __A23_NET_237, GND, __A23_NET_238, CCH11, __A23_NET_237, RCH11_n, __A23_NET_238, CH1114, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23052(__A23_NET_241, CHWL16_n, WCH11_n, __A23_NET_242, __A23_NET_241, __A23_NET_240, GND, __A23_NET_242, CCH11, __A23_NET_240, RCH11_n, __A23_NET_242, CH1116, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23053(__A23_NET_230, CHWL16_n, WCH12_n, __A23_NET_232, __A23_NET_230, __A23_NET_231, GND, __A23_NET_232, CCH12, __A23_NET_231, RCH12_n, __A23_NET_232, CH1216, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0) U23054(__A23_NET_232, __A23_2__ISSTDC,  ,  , __A23_NET_233, ALTEST, GND, __A23_1__P04A, P04_n, __A23_1__PIPSAM_n, __A23_1__PIPSAM, __A23_1__PIPAXp_n, PIPAXp, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23055(__A23_NET_229, CHWL16_n, WCH13_n, T6ON_n, __A23_NET_229, __A23_NET_228, GND, RCH13_n, T6ON_n, CH1316, CHWL10_n, WCH13_n, __A23_NET_234, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23056(__A23_NET_233, __A23_NET_234, __A23_NET_235, __A23_NET_235, __A23_NET_233, CCH13, GND, RCH13_n, __A23_NET_233, CH1310, __A23_1__PIPSAM_n, __A23_1__PIPAXp_n, __A23_1__PIPGXp, VCC, SIM_RST, SIM_CLK);
    U74HC27 U23057(PIPPLS_n, SB2_n,  ,  ,  ,  , GND,  ,  ,  ,  , __A23_1__PIPSAM, __A23_1__P04A, VCC, SIM_RST, SIM_CLK);
    U74HC04 U23058(PIPAXm, __A23_1__PIPAXm_n, PIPAYp, __A23_1__PIPAYp_n, PIPAYm, __A23_1__PIPAYm_n, GND, __A23_1__PIPAZp_n, PIPAZp, __A23_1__PIPAZm_n, PIPAZm,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U23059(__A23_1__PIPGXm, __A23_1__PIPSAM_n, __A23_1__PIPAXm_n, __A23_1__PIPGYp, __A23_1__PIPSAM_n, __A23_1__PIPAYp_n, GND, __A23_1__PIPSAM_n, __A23_1__PIPAYm_n, __A23_1__PIPGYm, __A23_1__PIPSAM_n, __A23_1__PIPAZp_n, __A23_1__PIPGZp, VCC, SIM_RST, SIM_CLK);
    U74HC02 U23060(__A23_1__PIPGZm, __A23_1__PIPSAM_n, __A23_1__PIPAZm_n,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
endmodule