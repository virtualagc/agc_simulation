`include "components/agc_parts.v"

module timer(VCC, GND, SIM_RST, CLOCK, PHS2, PHS2_n, PHS4, PHS4_n, RT, CT, CT_n, WT, WT_n, STOP, OVFSTB_n);
    input wire SIM_RST;
    wire ODDSET_n;
    wire NET_31;
    wire __cdiv2_c;
    wire __cdiv1_b;
    output wire CT_n;
    wire __cdiv1_d;
    output wire PHS2;
    input wire GND;
    wire __cdiv2_b;
    wire __oddset;
    wire __ovfstb_r5;
    wire RINGB_n;
    wire NET_24;
    output wire CT;
    wire NET_32;
    wire __cdiv2_d;
    wire __cdiv1_a;
    wire NET_26;
    wire __cdiv2_fs_n;
    input wire CLOCK;
    wire __cdiv2_a;
    output wire RT;
    wire __cdiv2_fs;
    output wire OVFSTB_n;
    output wire WT_n;
    wire RINGA_n;
    input wire STOP;
    wire __ovfstb_r2;
    output wire PHS4_n;
    output wire PHS4;
    wire __ovfstb_r1;
    input wire VCC;
    wire TT_n;
    wire EVNSET_n;
    wire __ovfstb_r3;
    output wire WT;
    wire __ovfstb_r6;
    output wire PHS2_n;
    wire EVNSET;
    wire __ovfstb_r4;

    U74HC04 U3(__cdiv1_d, NET_26, PHS2, PHS2_n, PHS4, PHS4_n, GND, NET_24, __cdiv1_b, CT, NET_24, CT_n, CT, VCC, SIM_RST);
    U74HC02 #(0, 1, 0, 0) U1(__cdiv1_d, NET_32, __cdiv1_b, NET_32, __cdiv1_b, NET_31, GND, NET_32, __cdiv1_a, NET_31, __cdiv1_a, NET_31, PHS2, VCC, SIM_RST);
    U74HC02 U6(__cdiv2_d, __cdiv2_fs_n, __cdiv2_b, __cdiv2_c, __cdiv2_a, __cdiv2_fs, GND, __cdiv2_b, __cdiv2_fs, __cdiv2_fs_n, __cdiv2_fs_n, __cdiv2_a, __cdiv2_fs, VCC, SIM_RST);
    U74HC04 U5(NET_32, WT, WT, WT_n, WT, TT_n, GND, __ovfstb_r5, __ovfstb_r4, __ovfstb_r6, __ovfstb_r5, OVFSTB_n, __ovfstb_r2, VCC, SIM_RST);
    U74HC04 U8(__cdiv2_d, RINGA_n, __oddset, ODDSET_n, __cdiv2_c, RINGB_n, GND, EVNSET, RINGB_n, EVNSET_n, EVNSET, RT, __cdiv1_a, VCC, SIM_RST);
    wire U4_8_NC;
    wire U4_9_NC;
    wire U4_10_NC;
    wire U4_11_NC;
    wire U4_12_NC;
    wire U4_13_NC;
    U74HC02 U4(PHS4, NET_26, __cdiv1_a, __oddset, STOP, RINGA_n, GND, U4_8_NC, U4_9_NC, U4_10_NC, U4_11_NC, U4_12_NC, U4_13_NC, VCC, SIM_RST);
    U74HC02 U9(__ovfstb_r1, CT_n, __ovfstb_r2, __ovfstb_r2, __ovfstb_r6, __ovfstb_r1, GND, __ovfstb_r4, __ovfstb_r2, __ovfstb_r3, __ovfstb_r3, __ovfstb_r1, __ovfstb_r4, VCC, SIM_RST);
    wire U2_8_NC;
    wire U2_9_NC;
    wire U2_10_NC;
    wire U2_11_NC;
    U74HC27 #(0, 1, 0) U2(__cdiv1_d, CLOCK, __cdiv1_b, CLOCK, PHS2, __cdiv1_a, GND, U2_8_NC, U2_9_NC, U2_10_NC, U2_11_NC, __cdiv1_b, __cdiv1_a, VCC, SIM_RST);
    wire U7_8_NC;
    wire U7_9_NC;
    wire U7_10_NC;
    wire U7_11_NC;
    U74HC27 #(0, 1, 0) U7(__cdiv2_d, NET_26, __cdiv2_b, NET_26, __cdiv2_c, __cdiv2_a, GND, U7_8_NC, U7_9_NC, U7_10_NC, U7_11_NC, __cdiv2_b, __cdiv2_a, VCC, SIM_RST);
endmodule