`include "components/agc_parts.v"

module scaler(VCC, GND, SIM_RST, FS01_n, RCHAT_n, RCHBT_n);
    input wire SIM_RST;
    wire __A01_2__CHBT11;
    wire __A01_1__scaler_s3__FS_n;
    wire __A01_1__F02A;
    wire NET_197;
    wire __A01_1__CHAT07;
    wire NET_209;
    wire __A01_1__CHAT10;
    wire __A01_1__FS12;
    wire __A01_2__FS25;
    wire __A01_1__FS15;
    wire __A01_1__F11A;
    wire NET_187;
    wire __A01_2__F30B;
    wire NET_177;
    wire NET_195;
    wire __A01_1__F06B;
    wire __A01_1__FS08;
    wire __A01_1__scaler_s7__FS_n;
    wire __A01_2__F19A;
    wire __A01_1__scaler_s16__FS_n;
    wire __A01_2__F18B;
    wire NET_184;
    wire __A01_1__F09A;
    wire __A01_2__scaler_s23__FS_n;
    wire __A01_1__FS06;
    wire __A01_2__FS22;
    wire __A01_2__F29B;
    wire NET_221;
    wire NET_203;
    wire NET_196;
    wire __A01_2__CHBT09;
    wire __A01_2__CHBT08;
    wire NET_230;
    wire __A01_1__F04B;
    wire __A01_1__F07B;
    wire __A01_2__CHBT05;
    wire NET_192;
    wire __A01_1__FS03;
    wire __A01_1__scaler_s8__FS_n;
    wire __A01_1__F02B;
    wire __A01_2__scaler_s29__FS_n;
    wire NET_190;
    wire NET_193;
    wire NET_216;
    wire __A01_2__CHBT07;
    wire __A01_2__FS26;
    wire __A01_2__CHBT02;
    wire NET_185;
    wire NET_155;
    wire __A01_2__CHBT04;
    wire NET_172;
    wire __A01_2__F20A;
    wire __A01_1__scaler_s9__FS_n;
    wire NET_225;
    wire __A01_1__FS13;
    wire __A01_1__CHAT06;
    wire NET_212;
    wire __A01_1__F16B;
    wire __A01_2__scaler_s19__FS_n;
    wire __A01_2__F31B;
    input wire GND;
    wire __A01_1__FS02;
    wire __A01_1__scaler_s2__FS_n;
    wire __A01_2__CHAT14;
    wire __A01_2__F32B;
    wire __A01_1__F17B;
    wire __A01_2__CHBT14;
    wire NET_180;
    wire NET_170;
    wire __A01_2__FS28;
    wire __A01_2__scaler_s33__FS_n;
    wire NET_171;
    wire __A01_1__F13B;
    wire __A01_2__F23A;
    wire __A01_2__F19B;
    wire __A01_1__CHAT08;
    wire NET_198;
    wire __A01_1__scaler_s15__FS_n;
    wire __A01_2__F22A;
    wire __A01_1__F09B;
    wire __A01_2__CHBT13;
    input wire VCC;
    wire __A01_2__FS27;
    wire NET_179;
    wire __A01_2__FS32;
    wire NET_174;
    wire __A01_1__scaler_s11__FS_n;
    wire __A01_2__CHBT01;
    wire __A01_1__FS16;
    wire __A01_1__F03A;
    wire __A01_1__F10A;
    wire __A01_2__scaler_s21__FS_n;
    wire __A01_2__F24B;
    wire NET_226;
    wire __A01_1__CHAT11;
    wire __A01_2__FS18;
    wire __A01_2__FS33;
    wire NET_223;
    wire __A01_1__scaler_s12__FS_n;
    wire __A01_1__F05A;
    wire __A01_1__FS11;
    wire NET_219;
    wire __A01_1__FS07;
    wire __A01_2__F22B;
    wire __A01_2__FS20;
    wire NET_173;
    wire NET_200;
    wire __A01_2__F21A;
    wire __A01_2__scaler_s26__FS_n;
    wire NET_189;
    wire __A01_2__F21B;
    wire __A01_2__F33A;
    wire NET_186;
    wire __A01_1__FS14;
    wire __A01_1__F15A;
    wire __A01_1__F03B;
    wire __A01_1__F17A;
    wire __A01_2__F26B;
    wire __A01_2__F25A;
    wire NET_194;
    wire __A01_1__FS03A;
    wire __A01_2__F30A;
    wire __A01_1__FS05;
    wire __A01_1__CHAT12;
    wire NET_201;
    wire __A01_1__F08A;
    wire __A01_1__FS04A;
    wire __A01_1__CHAT03;
    wire __A01_2__F28A;
    wire NET_143;
    wire __A01_1__FS09;
    wire NET_182;
    wire __A01_2__FS29;
    wire __A01_1__F04A;
    wire __A01_2__CHBT10;
    wire NET_207;
    wire NET_217;
    wire __A01_1__FS10;
    wire NET_181;
    wire __A01_1__F08B;
    wire __A01_2__CHBT06;
    wire __A01_1__FS02A;
    wire __A01_1__FS05A;
    wire NET_175;
    wire __A01_1__CHAT01;
    wire NET_211;
    wire __A01_1__F13A;
    wire __A01_2__FS24;
    wire __A01_1__F14B;
    wire NET_191;
    wire __A01_2__scaler_s32__FS_n;
    wire __A01_2__FS19;
    wire __A01_2__F27A;
    wire __A01_2__F24A;
    wire NET_228;
    wire __A01_1__CHAT02;
    wire __A01_1__F10B;
    wire __A01_1__scaler_s5__FS_n;
    wire __A01_1__CHAT04;
    wire __A01_2__F33B;
    wire __A01_1__scaler_s6__FS_n;
    wire NET_215;
    wire NET_178;
    wire NET_210;
    wire NET_206;
    wire NET_227;
    wire __A01_2__F28B;
    wire NET_229;
    wire __A01_2__F32A;
    wire __A01_2__CHAT13;
    wire __A01_1__F16A;
    wire NET_205;
    wire __A01_2__scaler_s30__FS_n;
    wire __A01_2__F18A;
    wire __A01_2__CHBT12;
    wire __A01_1__FS04;
    wire NET_218;
    wire __A01_1__CHAT09;
    wire __A01_1__F07A;
    input wire FS01_n;
    wire __A01_1__scaler_s10__FS_n;
    wire NET_224;
    wire __A01_1__scaler_s17__FS_n;
    wire NET_213;
    wire NET_204;
    wire NET_214;
    wire __A01_2__scaler_s20__FS_n;
    wire __A01_2__F25B;
    wire __A01_2__scaler_s18__FS_n;
    wire __A01_2__F26A;
    wire __A01_2__scaler_s22__FS_n;
    wire __A01_2__scaler_s27__FS_n;
    wire __A01_2__scaler_s24__FS_n;
    wire NET_188;
    wire NET_231;
    wire __A01_1__F15B;
    wire __A01_2__F23B;
    wire NET_183;
    wire __A01_2__FS30;
    wire __A01_1__F14A;
    input wire RCHBT_n;
    wire __A01_2__F29A;
    wire NET_222;
    wire __A01_1__scaler_s14__FS_n;
    wire __A01_2__FS23;
    wire __A01_2__F27B;
    wire __A01_2__scaler_s28__FS_n;
    input wire RCHAT_n;
    wire NET_208;
    wire __A01_2__FS21;
    wire __A01_1__F06A;
    wire NET_176;
    wire __A01_1__CHAT05;
    wire __A01_1__FS17;
    wire __A01_2__scaler_s31__FS_n;
    wire __A01_1__scaler_s13__FS_n;
    wire __A01_1__F11B;
    wire NET_169;
    wire __A01_1__F12B;
    wire NET_199;
    wire __A01_2__F20B;
    wire NET_202;
    wire __A01_2__CHBT03;
    wire __A01_2__FS31;
    wire __A01_2__scaler_s25__FS_n;
    wire NET_220;
    wire __A01_1__F12A;
    wire __A01_1__F05B;
    wire __A01_1__scaler_s4__FS_n;
    wire NET_168;
    wire __A01_2__F31A;

    U74HC02 #(0, 0, 1, 0) U1034(__A01_2__F19A, __A01_2__scaler_s19__FS_n, NET_203, __A01_2__F19B, NET_202, __A01_2__FS19, GND, NET_203, __A01_2__FS19, __A01_2__scaler_s19__FS_n, __A01_2__scaler_s19__FS_n, NET_202, __A01_2__FS19, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1011(__A01_1__F08A, __A01_1__scaler_s8__FS_n, NET_181, __A01_1__F08B, NET_180, __A01_1__FS08, GND, NET_181, __A01_1__FS08, __A01_1__scaler_s8__FS_n, __A01_1__scaler_s8__FS_n, NET_180, __A01_1__FS08, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1039(__A01_2__F22A, __A01_2__scaler_s22__FS_n, NET_209, __A01_2__F22B, NET_208, __A01_2__FS22, GND, NET_209, __A01_2__FS22, __A01_2__scaler_s22__FS_n, __A01_2__scaler_s22__FS_n, NET_208, __A01_2__FS22, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1003(__A01_1__F03A, __A01_1__scaler_s3__FS_n, NET_171, __A01_1__F03B, NET_170, __A01_1__FS03, GND, NET_171, __A01_1__FS03, __A01_1__scaler_s3__FS_n, __A01_1__scaler_s3__FS_n, NET_170, __A01_1__FS03, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1023(__A01_1__F15A, __A01_1__scaler_s15__FS_n, NET_195, __A01_1__F15B, NET_194, __A01_1__FS15, GND, NET_195, __A01_1__FS15, __A01_1__scaler_s15__FS_n, __A01_1__scaler_s15__FS_n, NET_194, __A01_1__FS15, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1006(__A01_1__F05A, __A01_1__scaler_s5__FS_n, NET_174, __A01_1__F05B, NET_175, __A01_1__FS05, GND, NET_174, __A01_1__FS05, __A01_1__scaler_s5__FS_n, __A01_1__scaler_s5__FS_n, NET_175, __A01_1__FS05, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1009(NET_176, __A01_1__F05A, __A01_1__F07A, __A01_1__F06A, NET_178, NET_179, GND, NET_178, NET_179, __A01_1__F06A, __A01_1__F07B, NET_177, __A01_1__F06B, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1017(__A01_1__F11A, __A01_1__F10A, NET_187, __A01_1__F10A, __A01_1__F11B, NET_186, GND, NET_188, __A01_1__F12A, __A01_1__F11A, NET_189, NET_187, NET_186, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1054(__A01_2__F31A, __A01_2__scaler_s31__FS_n, NET_227, __A01_2__F31B, NET_226, __A01_2__FS31, GND, NET_227, __A01_2__FS31, __A01_2__scaler_s31__FS_n, __A01_2__scaler_s31__FS_n, NET_226, __A01_2__FS31, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1057(__A01_2__F33A, __A01_2__scaler_s33__FS_n, NET_231, __A01_2__F33B, NET_230, __A01_2__FS33, GND, NET_231, __A01_2__FS33, __A01_2__scaler_s33__FS_n, __A01_2__scaler_s33__FS_n, NET_230, __A01_2__FS33, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1012(__A01_1__F08A, __A01_1__F07A, NET_181, __A01_1__F07A, __A01_1__F08B, NET_180, GND, NET_183, __A01_1__F09A, __A01_1__F08A, NET_182, NET_181, NET_180, VCC, SIM_RST);
    U74HC02 U1062(__A01_2__CHBT11, RCHBT_n, __A01_2__scaler_s30__FS_n, __A01_2__CHBT12, NET_155, __A01_2__scaler_s31__FS_n, GND, RCHBT_n, __A01_2__scaler_s32__FS_n, __A01_2__CHBT13, RCHBT_n, __A01_2__scaler_s33__FS_n, __A01_2__CHBT14, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1036(__A01_2__F20A, __A01_2__scaler_s20__FS_n, NET_205, __A01_2__F20B, NET_204, __A01_2__FS20, GND, NET_205, __A01_2__FS20, __A01_2__scaler_s20__FS_n, __A01_2__scaler_s20__FS_n, NET_204, __A01_2__FS20, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1020(__A01_1__F13A, __A01_1__scaler_s13__FS_n, NET_191, __A01_1__F13B, NET_190, __A01_1__FS13, GND, NET_191, __A01_1__FS13, __A01_1__scaler_s13__FS_n, __A01_1__scaler_s13__FS_n, NET_190, __A01_1__FS13, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1040(NET_209, __A01_2__F21A, __A01_2__F23A, __A01_2__F22A, NET_210, NET_211, GND, NET_210, NET_211, __A01_2__F22A, __A01_2__F23B, NET_208, __A01_2__F22B, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1041(__A01_2__F23A, __A01_2__scaler_s23__FS_n, NET_211, __A01_2__F23B, NET_210, __A01_2__FS23, GND, NET_211, __A01_2__FS23, __A01_2__scaler_s23__FS_n, __A01_2__scaler_s23__FS_n, NET_210, __A01_2__FS23, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1052(__A01_2__F30A, __A01_2__scaler_s30__FS_n, NET_225, __A01_2__F30B, NET_224, __A01_2__FS30, GND, NET_225, __A01_2__FS30, __A01_2__scaler_s30__FS_n, __A01_2__scaler_s30__FS_n, NET_224, __A01_2__FS30, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1010(__A01_1__F07A, __A01_1__scaler_s7__FS_n, NET_179, __A01_1__F07B, NET_178, __A01_1__FS07, GND, NET_179, __A01_1__FS07, __A01_1__scaler_s7__FS_n, __A01_1__scaler_s7__FS_n, NET_178, __A01_1__FS07, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1025(__A01_1__F16A, __A01_1__scaler_s16__FS_n, NET_196, __A01_1__F16B, NET_197, __A01_1__FS16, GND, NET_196, __A01_1__FS16, __A01_1__scaler_s16__FS_n, __A01_1__scaler_s16__FS_n, NET_197, __A01_1__FS16, VCC, SIM_RST);
    U74HC02 U1029(__A01_1__CHAT01, RCHAT_n, __A01_1__scaler_s6__FS_n, __A01_1__CHAT02, RCHAT_n, __A01_1__scaler_s7__FS_n, GND, RCHAT_n, __A01_1__scaler_s8__FS_n, __A01_1__CHAT03, RCHAT_n, __A01_1__scaler_s9__FS_n, __A01_1__CHAT04, VCC, SIM_RST);
    U74HC02 U1060(__A01_2__CHBT03, RCHBT_n, __A01_2__scaler_s22__FS_n, __A01_2__CHBT04, RCHBT_n, __A01_2__scaler_s23__FS_n, GND, RCHBT_n, __A01_2__scaler_s24__FS_n, __A01_2__CHBT05, RCHBT_n, __A01_2__scaler_s25__FS_n, __A01_2__CHBT06, VCC, SIM_RST);
    U74HC02 U1059(__A01_2__CHAT13, RCHAT_n, __A01_2__scaler_s18__FS_n, __A01_2__CHAT14, RCHAT_n, __A01_2__scaler_s19__FS_n, GND, RCHBT_n, __A01_2__scaler_s20__FS_n, __A01_2__CHBT01, RCHBT_n, __A01_2__scaler_s21__FS_n, __A01_2__CHBT02, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1026(__A01_1__F17A, __A01_1__scaler_s17__FS_n, NET_199, __A01_1__F17B, NET_198, __A01_1__FS17, GND, NET_199, __A01_1__FS17, __A01_1__scaler_s17__FS_n, __A01_1__scaler_s17__FS_n, NET_198, __A01_1__FS17, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1001(__A01_1__F02A, __A01_1__scaler_s2__FS_n, NET_169, __A01_1__F02B, NET_168, __A01_1__FS02, GND, NET_169, __A01_1__FS02, __A01_1__scaler_s2__FS_n, __A01_1__scaler_s2__FS_n, NET_168, __A01_1__FS02, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1043(__A01_2__F24A, __A01_2__F23A, NET_213, __A01_2__F23A, __A01_2__F24B, NET_212, GND, NET_215, __A01_2__F25A, __A01_2__F24A, NET_214, NET_213, NET_212, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1035(NET_203, __A01_2__F18A, __A01_2__F20A, __A01_2__F19A, NET_204, NET_205, GND, NET_204, NET_205, __A01_2__F19A, __A01_2__F20B, NET_202, __A01_2__F19B, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1022(__A01_1__F14A, __A01_1__F13A, NET_193, __A01_1__F13A, __A01_1__F14B, NET_192, GND, NET_195, __A01_1__F15A, __A01_1__F14A, NET_194, NET_193, NET_192, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1056(__A01_2__F32A, __A01_2__scaler_s32__FS_n, NET_229, __A01_2__F32B, NET_228, __A01_2__FS32, GND, NET_229, __A01_2__FS32, __A01_2__scaler_s32__FS_n, __A01_2__scaler_s32__FS_n, NET_228, __A01_2__FS32, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1024(NET_195, __A01_1__F14A, __A01_1__F16A, __A01_1__F15A, NET_197, NET_196, GND, NET_197, NET_196, __A01_1__F15A, __A01_1__F16B, NET_194, __A01_1__F15B, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1055(NET_227, __A01_2__F30A, __A01_2__F32A, __A01_2__F31A, NET_228, NET_229, GND, NET_228, NET_229, __A01_2__F31A, __A01_2__F32B, NET_226, __A01_2__F31B, VCC, SIM_RST);
    wire U1058_8_NC;
    wire U1058_9_NC;
    wire U1058_10_NC;
    wire U1058_11_NC;
    U74HC27 #(0, 1, 0) U1058(__A01_2__F33A, __A01_2__F32A, NET_231, __A01_2__F32A, __A01_2__F33B, NET_230, GND, U1058_8_NC, U1058_9_NC, U1058_10_NC, U1058_11_NC, NET_231, NET_230, VCC, SIM_RST);
    U74HC02 U1030(__A01_1__CHAT05, RCHAT_n, __A01_1__scaler_s10__FS_n, __A01_1__CHAT06, RCHAT_n, __A01_1__scaler_s11__FS_n, GND, RCHAT_n, __A01_1__scaler_s12__FS_n, __A01_1__CHAT07, RCHAT_n, __A01_1__scaler_s13__FS_n, __A01_1__CHAT08, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1002(__A01_1__F02A, FS01_n, NET_169, FS01_n, __A01_1__F02B, NET_168, GND, NET_171, __A01_1__F03A, __A01_1__F02A, NET_170, NET_169, NET_168, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1019(NET_188, __A01_1__F11A, __A01_1__F13A, __A01_1__F12A, NET_190, NET_191, GND, NET_190, NET_191, __A01_1__F12A, __A01_1__F13B, NET_189, __A01_1__F12B, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1016(__A01_1__F11A, __A01_1__scaler_s11__FS_n, NET_187, __A01_1__F11B, NET_186, __A01_1__FS11, GND, NET_187, __A01_1__FS11, __A01_1__scaler_s11__FS_n, __A01_1__scaler_s11__FS_n, NET_186, __A01_1__FS11, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1046(__A01_2__F26A, __A01_2__scaler_s26__FS_n, NET_217, __A01_2__F26B, NET_216, __A01_2__FS26, GND, NET_217, __A01_2__FS26, __A01_2__scaler_s26__FS_n, __A01_2__scaler_s26__FS_n, NET_216, __A01_2__FS26, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1013(__A01_1__F09A, __A01_1__scaler_s9__FS_n, NET_183, __A01_1__F09B, NET_182, __A01_1__FS09, GND, NET_183, __A01_1__FS09, __A01_1__scaler_s9__FS_n, __A01_1__scaler_s9__FS_n, NET_182, __A01_1__FS09, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1004(NET_171, __A01_1__F02A, __A01_1__F04A, __A01_1__F03A, NET_172, NET_173, GND, NET_172, NET_173, __A01_1__F03A, __A01_1__F04B, NET_170, __A01_1__F03B, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1005(__A01_1__F04A, __A01_1__scaler_s4__FS_n, NET_173, __A01_1__F04B, NET_172, __A01_1__FS04, GND, NET_173, __A01_1__FS04, __A01_1__scaler_s4__FS_n, __A01_1__scaler_s4__FS_n, NET_172, __A01_1__FS04, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1038(__A01_2__F21A, __A01_2__F20A, NET_207, __A01_2__F20A, __A01_2__F21B, NET_206, GND, NET_209, __A01_2__F22A, __A01_2__F21A, NET_208, NET_207, NET_206, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1008(__A01_1__F06A, __A01_1__scaler_s6__FS_n, NET_176, __A01_1__F06B, NET_177, __A01_1__FS06, GND, NET_176, __A01_1__FS06, __A01_1__scaler_s6__FS_n, __A01_1__scaler_s6__FS_n, NET_177, __A01_1__FS06, VCC, SIM_RST);
    wire U1027_8_NC;
    wire U1027_9_NC;
    wire U1027_10_NC;
    wire U1027_11_NC;
    U74HC27 #(0, 1, 0) U1027(__A01_1__F17A, __A01_1__F16A, NET_199, __A01_1__F16A, __A01_1__F17B, NET_198, GND, U1027_8_NC, U1027_9_NC, U1027_10_NC, U1027_11_NC, NET_199, NET_198, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1044(__A01_2__F25A, __A01_2__scaler_s25__FS_n, NET_215, __A01_2__F25B, NET_214, __A01_2__FS25, GND, NET_215, __A01_2__FS25, __A01_2__scaler_s25__FS_n, __A01_2__scaler_s25__FS_n, NET_214, __A01_2__FS25, VCC, SIM_RST);
    U74HC02 U1061(__A01_2__CHBT07, RCHBT_n, __A01_2__scaler_s26__FS_n, __A01_2__CHBT08, RCHBT_n, __A01_2__scaler_s27__FS_n, GND, RCHBT_n, __A01_2__scaler_s28__FS_n, __A01_2__CHBT09, RCHBT_n, __A01_2__scaler_s29__FS_n, __A01_2__CHBT10, VCC, SIM_RST);
    wire U1028_10_NC;
    wire U1028_11_NC;
    wire U1028_12_NC;
    wire U1028_13_NC;
    U74HC04 U1028(__A01_1__scaler_s2__FS_n, __A01_1__FS02A, __A01_1__scaler_s3__FS_n, __A01_1__FS03A, __A01_1__scaler_s4__FS_n, __A01_1__FS04A, GND, __A01_1__FS05A, __A01_1__scaler_s5__FS_n, U1028_10_NC, U1028_11_NC, U1028_12_NC, U1028_13_NC, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1015(__A01_1__F10A, __A01_1__scaler_s10__FS_n, NET_185, __A01_1__F10B, NET_184, __A01_1__FS10, GND, NET_185, __A01_1__FS10, __A01_1__scaler_s10__FS_n, __A01_1__scaler_s10__FS_n, NET_184, __A01_1__FS10, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1042(__A01_2__F24A, __A01_2__scaler_s24__FS_n, NET_213, __A01_2__F24B, NET_212, __A01_2__FS24, GND, NET_213, __A01_2__FS24, __A01_2__scaler_s24__FS_n, __A01_2__scaler_s24__FS_n, NET_212, __A01_2__FS24, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1033(__A01_2__F18A, __A01_1__F17A, NET_201, __A01_1__F17A, __A01_2__F18B, NET_200, GND, NET_203, __A01_2__F19A, __A01_2__F18A, NET_202, NET_201, NET_200, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1049(__A01_2__F28A, __A01_2__scaler_s28__FS_n, NET_221, __A01_2__F28B, NET_220, __A01_2__FS28, GND, NET_221, __A01_2__FS28, __A01_2__scaler_s28__FS_n, __A01_2__scaler_s28__FS_n, NET_220, __A01_2__FS28, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1007(__A01_1__F05A, __A01_1__F04A, NET_174, __A01_1__F04A, __A01_1__F05B, NET_175, GND, NET_176, __A01_1__F06A, __A01_1__F05A, NET_177, NET_174, NET_175, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1037(__A01_2__F21A, __A01_2__scaler_s21__FS_n, NET_207, __A01_2__F21B, NET_206, __A01_2__FS21, GND, NET_207, __A01_2__FS21, __A01_2__scaler_s21__FS_n, __A01_2__scaler_s21__FS_n, NET_206, __A01_2__FS21, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1032(__A01_2__F18A, __A01_2__scaler_s18__FS_n, NET_201, __A01_2__F18B, NET_200, __A01_2__FS18, GND, NET_201, __A01_2__FS18, __A01_2__scaler_s18__FS_n, __A01_2__scaler_s18__FS_n, NET_200, __A01_2__FS18, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1021(__A01_1__F14A, __A01_1__scaler_s14__FS_n, NET_193, __A01_1__F14B, NET_192, __A01_1__FS14, GND, NET_193, __A01_1__FS14, __A01_1__scaler_s14__FS_n, __A01_1__scaler_s14__FS_n, NET_192, __A01_1__FS14, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1048(__A01_2__F27A, __A01_2__F26A, NET_219, __A01_2__F26A, __A01_2__F27B, NET_218, GND, NET_221, __A01_2__F28A, __A01_2__F27A, NET_220, NET_219, NET_218, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1051(__A01_2__F29A, __A01_2__scaler_s29__FS_n, NET_223, __A01_2__F29B, NET_222, __A01_2__FS29, GND, NET_223, __A01_2__FS29, __A01_2__scaler_s29__FS_n, __A01_2__scaler_s29__FS_n, NET_222, __A01_2__FS29, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1047(__A01_2__F27A, __A01_2__scaler_s27__FS_n, NET_219, __A01_2__F27B, NET_218, __A01_2__FS27, GND, NET_219, __A01_2__FS27, __A01_2__scaler_s27__FS_n, __A01_2__scaler_s27__FS_n, NET_218, __A01_2__FS27, VCC, SIM_RST);
    U74HC02 U1031(__A01_1__CHAT09, RCHAT_n, __A01_1__scaler_s14__FS_n, __A01_1__CHAT10, NET_143, __A01_1__scaler_s15__FS_n, GND, RCHAT_n, __A01_1__scaler_s16__FS_n, __A01_1__CHAT11, RCHAT_n, __A01_1__scaler_s17__FS_n, __A01_1__CHAT12, VCC, SIM_RST);
    U74HC02 #(0, 0, 1, 0) U1018(__A01_1__F12A, __A01_1__scaler_s12__FS_n, NET_188, __A01_1__F12B, NET_189, __A01_1__FS12, GND, NET_188, __A01_1__FS12, __A01_1__scaler_s12__FS_n, __A01_1__scaler_s12__FS_n, NET_189, __A01_1__FS12, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1050(NET_221, __A01_2__F27A, __A01_2__F29A, __A01_2__F28A, NET_222, NET_223, GND, NET_222, NET_223, __A01_2__F28A, __A01_2__F29B, NET_220, __A01_2__F28B, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1014(NET_183, __A01_1__F08A, __A01_1__F10A, __A01_1__F09A, NET_184, NET_185, GND, NET_184, NET_185, __A01_1__F09A, __A01_1__F10B, NET_182, __A01_1__F09B, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1045(NET_215, __A01_2__F24A, __A01_2__F26A, __A01_2__F25A, NET_216, NET_217, GND, NET_216, NET_217, __A01_2__F25A, __A01_2__F26B, NET_214, __A01_2__F25B, VCC, SIM_RST);
    U74HC27 #(0, 1, 0) U1053(__A01_2__F30A, __A01_2__F29A, NET_225, __A01_2__F29A, __A01_2__F30B, NET_224, GND, NET_227, __A01_2__F31A, __A01_2__F30A, NET_226, NET_225, NET_224, VCC, SIM_RST);
endmodule