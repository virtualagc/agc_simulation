`timescale 1ns/1ps
`default_nettype none

module fpga_agc(VCC, GND, SIM_RST, SIM_CLK, ALTEST, BLKUPL_n, BMGXM, BMGXP, BMGYM, BMGYP, BMGZM, BMGZP, CAURST, CCH13, CCH14, CCH34, CCH35, CDUFAL, CDUSTB_n, CDUXD, CDUXM, CDUXP, CDUYD, CDUYM, CDUYP, CDUZD, CDUZM, CDUZP, CH01, CH02, CH03, CH04, CH05, CH06, CH07, CH0705, CH0706, CH0707, CH08, CH09, CH10, CH11, CH12, CH13, CH1309, CH1310, CH1316, CH14, CH1411, CH1412, CH1413, CH1414, CH1416, CH16, CHWL01_n, CHWL02_n, CHWL03_n, CHWL04_n, CHWL05_n, CHWL06_n, CHWL07_n, CHWL08_n, CHWL09_n, CHWL10_n, CHWL11_n, CHWL12_n, CHWL13_n, CHWL14_n, CHWL16_n, CLOCK, CTLSAT, DBLTEST, DKBSNC, DKEND, DKSTRT, E5, E6, E7_n, EPCS_DATA, FLASH, FLASH_n, FLTOUT, FREFUN, GATEX_n, GATEY_n, GATEZ_n, GCAPCL, GTONE, GTRST_n, GTSET, GTSET_n, GUIREL, HNDRPT, HOLFUN, IMUCAG, IMUFAL, IMUOPR, IN3008, IN3212, IN3213, IN3214, IN3216, IN3301, ISSTOR, LEMATT, LFTOFF, LRIN0, LRIN1, LRRLSC, LVDAGD, MAINRS, MAMU, MANmP, MANmR, MANmY, MANpP, MANpR, MANpY, MARK, MDT01, MDT02, MDT03, MDT04, MDT05, MDT06, MDT07, MDT08, MDT09, MDT10, MDT11, MDT12, MDT13, MDT14, MDT15, MDT16, MKEY1, MKEY2, MKEY3, MKEY4, MKEY5, MLDCH, MLOAD, MNHNC, MNHRPT, MNHSBF, MNIMmP, MNIMmR, MNIMmY, MNIMpP, MNIMpR, MNIMpY, MONPAR, MONWBK, MRDCH, MREAD, MRKREJ, MRKRST, MSTP, MSTRT, MTCSAI, NAVRST, NHALGA, NHVFAL, NKEY1, NKEY2, NKEY3, NKEY4, NKEY5, OPCDFL, OPMSW2, OPMSW3, OVNHRP, PCHGOF, PIPAFL, PIPPLS_n, PIPXM, PIPXP, PIPYM, PIPYP, PIPZM, PIPZP, RCH13_n, RCH14_n, RCH33_n, RCHAT_n, RCHBT_n, ROLGOF, RRIN0, RRIN1, RRPONA, RRRLSC, S4BSAB, SBYBUT, SCAFAL, SHAFTD, SHAFTM, SHAFTP, SIGNX, SIGNY, SIGNZ, SMSEPR, SPSRDY, STRPRS, STRT2, T6ON_n, TEMPIN, TEMPIN_n, TRANmX, TRANmY, TRANmZ, TRANpX, TRANpY, TRANpZ, TRNM, TRNP, TRST10, TRST9, TRUND, ULLTHR, UPL0, UPL1, UPRUPT, VFAIL, WCH13_n, WCH14_n, WCH34_n, WCH35_n, XLNK0, XLNK1, ZEROP, n2FSFAL, EPCS_ASDI, EPCS_CSN, EPCS_DCLK, MGOJAM, MT01, MT02, MT03, MT04, MT05, MT06, MT07, MT08, MT09, MT10, MT11, MT12);
    input wire VCC;
    input wire GND;
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire ALTEST;
    input wire BLKUPL_n;
    input wire BMGXM;
    input wire BMGXP;
    input wire BMGYM;
    input wire BMGYP;
    input wire BMGZM;
    input wire BMGZP;
    input wire CAURST;
    input wire CCH13;
    input wire CCH14;
    input wire CCH34;
    input wire CCH35;
    input wire CDUFAL;
    input wire CDUSTB_n;
    input wire CDUXD;
    input wire CDUXM;
    input wire CDUXP;
    input wire CDUYD;
    input wire CDUYM;
    input wire CDUYP;
    input wire CDUZD;
    input wire CDUZM;
    input wire CDUZP;
    input wire CH01;
    input wire CH02;
    input wire CH03;
    input wire CH04;
    input wire CH05;
    input wire CH06;
    input wire CH07;
    input wire CH0705;
    input wire CH0706;
    input wire CH0707;
    input wire CH08;
    input wire CH09;
    input wire CH10;
    input wire CH11;
    input wire CH12;
    input wire CH13;
    input wire CH1309;
    input wire CH1310;
    input wire CH1316;
    input wire CH14;
    input wire CH1411;
    input wire CH1412;
    input wire CH1413;
    input wire CH1414;
    input wire CH1416;
    input wire CH16;
    input wire CHWL01_n;
    input wire CHWL02_n;
    input wire CHWL03_n;
    input wire CHWL04_n;
    input wire CHWL05_n;
    input wire CHWL06_n;
    input wire CHWL07_n;
    input wire CHWL08_n;
    input wire CHWL09_n;
    input wire CHWL10_n;
    input wire CHWL11_n;
    input wire CHWL12_n;
    input wire CHWL13_n;
    input wire CHWL14_n;
    input wire CHWL16_n;
    input wire CLOCK;
    input wire CTLSAT;
    input wire DBLTEST;
    input wire DKBSNC;
    input wire DKEND;
    input wire DKSTRT;
    input wire E5;
    input wire E6;
    input wire E7_n;
    input wire EPCS_DATA;
    input wire FLASH;
    input wire FLASH_n;
    input wire FLTOUT;
    input wire FREFUN;
    input wire GATEX_n;
    input wire GATEY_n;
    input wire GATEZ_n;
    input wire GCAPCL;
    input wire GTONE;
    input wire GTRST_n;
    input wire GTSET;
    input wire GTSET_n;
    input wire GUIREL;
    input wire HNDRPT;
    input wire HOLFUN;
    input wire IMUCAG;
    input wire IMUFAL;
    input wire IMUOPR;
    input wire IN3008;
    input wire IN3212;
    input wire IN3213;
    input wire IN3214;
    input wire IN3216;
    input wire IN3301;
    input wire ISSTOR;
    input wire LEMATT;
    input wire LFTOFF;
    input wire LRIN0;
    input wire LRIN1;
    input wire LRRLSC;
    input wire LVDAGD;
    input wire MAINRS;
    input wire MAMU;
    input wire MANmP;
    input wire MANmR;
    input wire MANmY;
    input wire MANpP;
    input wire MANpR;
    input wire MANpY;
    input wire MARK;
    input wire MDT01;
    input wire MDT02;
    input wire MDT03;
    input wire MDT04;
    input wire MDT05;
    input wire MDT06;
    input wire MDT07;
    input wire MDT08;
    input wire MDT09;
    input wire MDT10;
    input wire MDT11;
    input wire MDT12;
    input wire MDT13;
    input wire MDT14;
    input wire MDT15;
    input wire MDT16;
    input wire MKEY1;
    input wire MKEY2;
    input wire MKEY3;
    input wire MKEY4;
    input wire MKEY5;
    input wire MLDCH;
    input wire MLOAD;
    input wire MNHNC;
    input wire MNHRPT;
    input wire MNHSBF;
    input wire MNIMmP;
    input wire MNIMmR;
    input wire MNIMmY;
    input wire MNIMpP;
    input wire MNIMpR;
    input wire MNIMpY;
    input wire MONPAR;
    input wire MONWBK;
    input wire MRDCH;
    input wire MREAD;
    input wire MRKREJ;
    input wire MRKRST;
    input wire MSTP;
    input wire MSTRT;
    input wire MTCSAI;
    input wire NAVRST;
    input wire NHALGA;
    input wire NHVFAL;
    input wire NKEY1;
    input wire NKEY2;
    input wire NKEY3;
    input wire NKEY4;
    input wire NKEY5;
    input wire OPCDFL;
    input wire OPMSW2;
    input wire OPMSW3;
    input wire OVNHRP;
    input wire PCHGOF;
    input wire PIPAFL;
    input wire PIPPLS_n;
    input wire PIPXM;
    input wire PIPXP;
    input wire PIPYM;
    input wire PIPYP;
    input wire PIPZM;
    input wire PIPZP;
    input wire RCH13_n;
    input wire RCH14_n;
    input wire RCH33_n;
    input wire RCHAT_n;
    input wire RCHBT_n;
    input wire ROLGOF;
    input wire RRIN0;
    input wire RRIN1;
    input wire RRPONA;
    input wire RRRLSC;
    input wire S4BSAB;
    input wire SBYBUT;
    input wire SCAFAL;
    input wire SHAFTD;
    input wire SHAFTM;
    input wire SHAFTP;
    input wire SIGNX;
    input wire SIGNY;
    input wire SIGNZ;
    input wire SMSEPR;
    input wire SPSRDY;
    input wire STRPRS;
    input wire STRT2;
    input wire T6ON_n;
    input wire TEMPIN;
    input wire TEMPIN_n;
    input wire TRANmX;
    input wire TRANmY;
    input wire TRANmZ;
    input wire TRANpX;
    input wire TRANpY;
    input wire TRANpZ;
    input wire TRNM;
    input wire TRNP;
    input wire TRST10;
    input wire TRST9;
    input wire TRUND;
    input wire ULLTHR;
    input wire UPL0;
    input wire UPL1;
    input wire UPRUPT;
    input wire VFAIL;
    input wire WCH13_n;
    input wire WCH14_n;
    input wire WCH34_n;
    input wire WCH35_n;
    input wire XLNK0;
    input wire XLNK1;
    input wire ZEROP;
    input wire n2FSFAL;
    output wire EPCS_ASDI;
    output wire EPCS_CSN;
    output wire EPCS_DCLK;
    output wire MGOJAM;
    output wire MT01;
    output wire MT02;
    output wire MT03;
    output wire MT04;
    output wire MT05;
    output wire MT06;
    output wire MT07;
    output wire MT08;
    output wire MT09;
    output wire MT10;
    output wire MT11;
    output wire MT12;
    wire A2XG_n;
    wand A2X_n;
    wire A2X_n_U5012_10;
    wire A2X_n_U5046_8;
    wire A2X_n_U6004_6;
    wire AD0;
    wire ADS0;
    wire AGCWAR;
    wire ALGA;
    wire ALTM;
    wire AUG0_n;
    wire B15X;
    wire BKTF_n;
    wire BMAGXM;
    wire BMAGXP;
    wire BMAGYM;
    wire BMAGYP;
    wire BMAGZM;
    wire BMAGZP;
    wire BR1;
    wire BR12B_n;
    wire BR1B2B;
    wire BR1B2B_n;
    wire BR1B2_n;
    wire BR1_n;
    wire BR2;
    wire BR2_n;
    wire BRDIF_n;
    wire BXVX;
    wire C24A;
    wire C25A;
    wire C26A;
    wire C27A;
    wire C30A;
    wire C31A;
    wire C32A;
    wire C32M;
    wire C32P;
    wire C33A;
    wire C33M;
    wire C33P;
    wire C34A;
    wire C34M;
    wire C34P;
    wire C35A;
    wire C35M;
    wire C35P;
    wire C36A;
    wire C36M;
    wire C36P;
    wire C37A;
    wire C37M;
    wire C37P;
    wire C40A;
    wire C40M;
    wire C40P;
    wire C41A;
    wire C41M;
    wire C41P;
    wire C45R;
    wire C50A;
    wire C51A;
    wire C52A;
    wire C53A;
    wire C54A;
    wire C55A;
    wire CA2_n;
    wire CA3_n;
    wire CA4_n;
    wire CA5_n;
    wire CA6_n;
    wire CAD1;
    wire CAD2;
    wire CAD3;
    wire CAD4;
    wire CAD5;
    wire CAD6;
    wire CAG;
    wire CBG;
    wire CCH11;
    wire CCH33;
    wire CCHG_n;
    wire CCS0;
    wire CCS0_n;
    wire CEBG;
    wire CFBG;
    wire CG13;
    wire CG23;
    wire CG26;
    wire CGG;
    wire CGMC;
    wire CH1213;
    wire CH1214;
    wire CH1301;
    wire CH1302;
    wire CH1303;
    wire CH1304;
    wire CH1305;
    wire CH1306;
    wire CH1307;
    wire CH1308;
    wire CH1311;
    wire CH1401;
    wire CH1402;
    wire CH1403;
    wire CH1404;
    wire CH1405;
    wire CH1406;
    wire CH1407;
    wire CH1408;
    wire CH1409;
    wire CH1410;
    wire CH1501;
    wire CH1502;
    wire CH1503;
    wire CH1504;
    wire CH3201;
    wire CH3202;
    wire CH3203;
    wire CH3204;
    wire CH3205;
    wire CH3206;
    wire CH3207;
    wire CH3208;
    wire CH3310;
    wire CH3312;
    wire CHINC;
    wire CHINC_n;
    wire CI01_n;
    wire CI05_n;
    wire CI09_n;
    wire CI13_n;
    wand CI_n;
    wire CI_n_U4061_12;
    wire CI_n_U5018_2;
    wire CI_n_U5046_10;
    wire CI_n_U6047_2;
    wire CLG1G;
    wire CLG2G;
    wire CLK;
    wire CLROPE;
    wire CLXC;
    wand CO06;
    wire CO06_U8041_2;
    wire CO06_U8050_2;
    wand CO10;
    wire CO10_U9041_2;
    wire CO10_U9050_2;
    wand CO14;
    wire CO14_U10041_2;
    wire CO14_U10050_2;
    wire CQG;
    wire CSG;
    wire CT;
    wire CTROR;
    wire CTROR_n;
    wire CT_n;
    wire CUG;
    wire CXB0_n;
    wire CXB1_n;
    wire CXB2_n;
    wire CXB3_n;
    wire CXB4_n;
    wire CXB5_n;
    wire CXB6_n;
    wire CXB7_n;
    wire CYL_n;
    wire CYR_n;
    wire CZG;
    wire DAS0;
    wire DAS0_n;
    wire DAS1;
    wire DAS1_n;
    wire DCA0;
    wire DCS0;
    wire DIM0_n;
    wire DINC;
    wire DINC_n;
    wire DIVSTG;
    wire DIV_n;
    wire DLKPLS;
    wire DRPRST;
    wire DV1;
    wire DV1376;
    wire DV1376_n;
    wire DV1_n;
    wire DV3764;
    wire DV376_n;
    wire DV4;
    wire DV4B1B;
    wire DV4_n;
    wire DVST;
    wire DXCH0;
    wire EAC_n;
    wire EB10;
    wire EB11_n;
    wire EB9;
    wire EDOP_n;
    wire EMSD;
    wire EXST0_n;
    wire EXST1_n;
    wire EXT;
    wire EXTPLS;
    wire F04A;
    wire F04B;
    wire F05A_n;
    wire F05B_n;
    wire F06B;
    wire F07A;
    wire F07B;
    wire F07B_n;
    wire F08B;
    wire F09A;
    wire F09B;
    wire F09B_n;
    wire F10A;
    wire F10A_n;
    wire F10B;
    wire F12B;
    wire F14B;
    wire F17A;
    wire F17B;
    wire F5ASB2_n;
    wire F5BSB2_n;
    wire FETCH0;
    wire FETCH0_n;
    wire FETCH1;
    wire FS01;
    wire FS01_n;
    wire FS05_n;
    wire FS07A;
    wire FS07_n;
    wire FS09;
    wire FS09_n;
    wire FS10;
    wire FS13;
    wire FS14;
    wire FUTEXT;
    wire G01;
    wire G01ED;
    wand G01_n;
    wire G01_n_U8013_6;
    wire G01_n_U8013_8;
    wire G02;
    wire G02ED;
    wire G03;
    wire G03ED;
    wire G04;
    wire G04ED;
    wire G05;
    wire G05ED;
    wand G05_n;
    wire G05_n_U9013_6;
    wire G05_n_U9013_8;
    wire G06;
    wire G06ED;
    wand G06_n;
    wire G06_n_U9028_10;
    wire G06_n_U9028_12;
    wire G07;
    wire G07ED;
    wand G07_n;
    wire G07_n_U9050_6;
    wire G07_n_U9050_8;
    wire G08;
    wire G09;
    wand G09_n;
    wire G09_n_U10013_6;
    wire G09_n_U10013_8;
    wire G10;
    wand G10_n;
    wire G10_n_U10028_10;
    wire G10_n_U10028_12;
    wire G11;
    wand G11_n;
    wire G11_n_U10050_6;
    wire G11_n_U10050_8;
    wire G12;
    wire G13;
    wand G13_n;
    wire G13_n_U11013_6;
    wire G13_n_U11013_8;
    wire G14;
    wand G14_n;
    wire G14_n_U11028_10;
    wire G14_n_U11028_12;
    wire G15;
    wand G15_n;
    wire G15_n_U11050_6;
    wire G15_n_U11050_8;
    wire G16;
    wire G16SW_n;
    wire G2LSG_n;
    wire GEM01;
    wire GEM02;
    wire GEM03;
    wire GEM04;
    wire GEM05;
    wire GEM06;
    wire GEM07;
    wire GEM08;
    wire GEM09;
    wire GEM10;
    wire GEM11;
    wire GEM12;
    wire GEM13;
    wire GEM14;
    wire GEM16;
    wire GEMP;
    wire GEQZRO_n;
    wire GINH;
    wire GNHNC;
    wire GOJ1;
    wire GOJ1_n;
    wire GOJAM;
    wire GOJAM_n;
    wire GYROD;
    wire HIMOD;
    wire IC1;
    wire IC10;
    wire IC10_n;
    wire IC11;
    wire IC11_n;
    wire IC12;
    wire IC12_n;
    wire IC13;
    wire IC14;
    wire IC15;
    wire IC15_n;
    wire IC16;
    wire IC16_n;
    wire IC17;
    wire IC2;
    wire IC2_n;
    wire IC3;
    wire IC4;
    wire IC5;
    wire IC5_n;
    wire IC6;
    wire IC7;
    wire IC8_n;
    wire IC9;
    wire IIP;
    wire IIP_n;
    wire IL01;
    wire IL02;
    wire IL03;
    wire IL04;
    wire IL05;
    wire IL06;
    wire IL07;
    wire INCR0;
    wire INCSET_n;
    wand INHPLS;
    wire INHPLS_U12016_10;
    wire INHPLS_U12016_12;
    wire INKL;
    wire INKL_n;
    wire INLNKM;
    wire INLNKP;
    wire INOTLD;
    wire INOUT;
    wire INOUT_n;
    wire KRPT;
    wire KYRPT1;
    wire KYRPT2;
    wand L01_n;
    wire L01_n_U8007_6;
    wand L02_n;
    wire L02_n_U8013_12;
    wand L04_n;
    wire L04_n_U8050_12;
    wand L08_n;
    wire L08_n_U9050_12;
    wand L12_n;
    wire L12_n_U10050_12;
    wand L15_n;
    wire L15_n_U11041_6;
    wand L16_n;
    wire L16_n_U11050_12;
    wire L16_n_U4063_8;
    wire L2GDG_n;
    wire L2GD_n;
    wire LOMOD;
    wire MASK0;
    wire MASK0_n;
    wire MCDU;
    wire MCRO_n;
    wire MINC;
    wire MKRPT;
    wire MONEX;
    wand MONEX_n;
    wire MONEX_n_U5005_2;
    wire MONEX_n_U6029_6;
    wire MONWT;
    wire MON_n;
    wire MONpCH;
    wire MOUT_n;
    wire MP0;
    wire MP0T10;
    wire MP0_n;
    wire MP1;
    wire MP1_n;
    wire MP3;
    wire MP3A;
    wire MP3_n;
    wire MSTPIT_n;
    wire MSTRTP;
    wire MSU0;
    wire MSU0_n;
    wire NDR100_n;
    wire NDX0_n;
    wire NDXX1_n;
    wire NEAC;
    wire NISQ;
    wire NISQL_n;
    wire OCTAD2;
    wire OCTAD3;
    wire OCTAD4;
    wire OCTAD5;
    wire OCTAD6;
    wire OSCALM;
    wire OTLNKM;
    wire OVF_n;
    wire P01;
    wire P01_n;
    wire P02;
    wire P02_n;
    wire P03;
    wire P03_n;
    wire P04;
    wire P04_n;
    wire P05;
    wire P05_n;
    wand PALE;
    wire PALE_U12027_2;
    wire PALE_U12027_4;
    wire PC15_n;
    wire PCDU;
    wire PHS2;
    wire PHS2_n;
    wire PHS3_n;
    wire PHS4;
    wire PHS4_n;
    wire PIFL_n;
    wire PINC;
    wire PONEX;
    wire POUT_n;
    wire PRINC;
    wire PSEUDO;
    wire PTWOX;
    wire Q2A;
    wire QC0_n;
    wire QC1_n;
    wire QC2_n;
    wire QC3_n;
    wire QXCH0_n;
    wire R15;
    wire R1C;
    wand R1C_n;
    wire R1C_n_U4063_10;
    wire R1C_n_U6029_12;
    wire R6;
    wire RAD;
    wire RADRG;
    wire RADRPT;
    wire RADRZ;
    wire RAG_n;
    wire RAND0;
    wand RA_n;
    wire RA_n_U4039_10;
    wire RA_n_U4045_8;
    wire RA_n_U5005_8;
    wire RA_n_U5024_4;
    wire RA_n_U5041_12;
    wire RB1;
    wire RB1F;
    wand RB1_n;
    wire RB1_n_U4063_6;
    wire RB1_n_U6029_10;
    wire RB2;
    wire RBBEG_n;
    wire RBHG_n;
    wire RBLG_n;
    wire RBSQ;
    wand RB_n;
    wire RB_n_U4039_2;
    wire RB_n_U4061_10;
    wire RB_n_U5005_6;
    wire RB_n_U5018_10;
    wire RB_n_U5051_2;
    wire RB_n_U6004_8;
    wire RB_n_U6037_8;
    wire RCG_n;
    wire RCH11_n;
    wire RCH_n;
    wand RC_n;
    wire RC_n_U4039_4;
    wire RC_n_U4061_8;
    wire RC_n_U5012_8;
    wire RC_n_U5024_10;
    wire RC_n_U5051_10;
    wire RC_n_U6047_6;
    wire RC_n_U6052_8;
    wire READ0;
    wire REBG_n;
    wand RELPLS;
    wire RELPLS_U12016_6;
    wire RELPLS_U12016_8;
    wire RESETA;
    wire RESETB;
    wire RESETC;
    wire RESETD;
    wire RFBG_n;
    wire RGG_n;
    wand RG_n;
    wire RG_n_U5012_6;
    wire RG_n_U5046_2;
    wire RG_n_U5046_4;
    wire RG_n_U5061_10;
    wire RG_n_U6014_8;
    wand RL01_n;
    wire RL01_n_U15039_12;
    wire RL01_n_U8007_10;
    wire RL01_n_U8007_12;
    wire RL01_n_U8007_4;
    wire RL01_n_U8013_4;
    wand RL02_n;
    wire RL02_n_U15039_10;
    wire RL02_n_U8013_10;
    wire RL02_n_U8028_2;
    wire RL02_n_U8028_6;
    wire RL02_n_U8028_8;
    wand RL03_n;
    wire RL03_n_U15039_4;
    wire RL03_n_U8041_10;
    wire RL03_n_U8041_12;
    wire RL03_n_U8041_4;
    wire RL03_n_U8050_4;
    wand RL04_n;
    wire RL04_n_U15039_6;
    wire RL04_n_U8050_10;
    wire RL04_n_U8063_2;
    wire RL04_n_U8063_6;
    wire RL04_n_U8063_8;
    wand RL05_n;
    wire RL05_n_U15039_8;
    wire RL05_n_U9007_10;
    wire RL05_n_U9007_12;
    wire RL05_n_U9007_4;
    wire RL05_n_U9013_4;
    wand RL06_n;
    wire RL06_n_U15016_6;
    wire RL06_n_U9013_10;
    wire RL06_n_U9028_2;
    wire RL06_n_U9028_6;
    wire RL06_n_U9028_8;
    wand RL09_n;
    wire RL09_n_U10007_10;
    wire RL09_n_U10007_12;
    wire RL09_n_U10007_4;
    wire RL09_n_U10013_4;
    wire RL09_n_U15016_4;
    wire RL10BB;
    wand RL10_n;
    wire RL10_n_U10013_10;
    wire RL10_n_U10028_2;
    wire RL10_n_U10028_6;
    wire RL10_n_U10028_8;
    wire RL10_n_U15016_2;
    wand RL11_n;
    wire RL11_n_U10041_10;
    wire RL11_n_U10041_12;
    wire RL11_n_U10041_4;
    wire RL11_n_U10050_4;
    wire RL11_n_U15004_12;
    wand RL12_n;
    wire RL12_n_U10050_10;
    wire RL12_n_U10063_2;
    wire RL12_n_U10063_6;
    wire RL12_n_U10063_8;
    wire RL12_n_U15004_10;
    wand RL13_n;
    wire RL13_n_U11007_10;
    wire RL13_n_U11007_12;
    wire RL13_n_U11007_4;
    wire RL13_n_U11013_4;
    wire RL13_n_U15004_8;
    wand RL14_n;
    wire RL14_n_U11013_10;
    wire RL14_n_U11028_2;
    wire RL14_n_U11028_6;
    wire RL14_n_U11028_8;
    wire RL14_n_U15004_6;
    wand RL15_n;
    wire RL15_n_U11041_10;
    wire RL15_n_U11041_12;
    wire RL15_n_U11041_4;
    wire RL15_n_U11050_4;
    wire RL15_n_U15004_4;
    wand RL16_n;
    wire RL16_n_U11050_10;
    wire RL16_n_U11063_2;
    wire RL16_n_U11063_6;
    wire RL16_n_U11063_8;
    wire RL16_n_U15004_2;
    wire RLG_n;
    wand RL_n;
    wire RL_n_U5005_12;
    wire RL_n_U5041_10;
    wire RNRADM;
    wire RNRADP;
    wire ROPER;
    wire ROPES;
    wire ROPET;
    wire ROR0;
    wand RPTSET;
    wire RPTSET_U3011_2;
    wire RPTSET_U3011_4;
    wire RPTSET_U3011_6;
    wire RPTSET_U6052_4;
    wire RQG_n;
    wire RQ_n;
    wire RRPA;
    wire RSCT;
    wire RSC_n;
    wire RSM3;
    wire RSM3_n;
    wire RSSB;
    wire RSTRT;
    wire RSTSTG;
    wire RT;
    wire RT_n;
    wire RUG_n;
    wire RULOG_n;
    wire RUPT0;
    wire RUPT1;
    wire RUPTOR_n;
    wire RUS_n;
    wand RU_n;
    wire RU_n_U5024_2;
    wire RU_n_U5061_4;
    wire RU_n_U5061_6;
    wire RU_n_U6014_12;
    wire RU_n_U6037_2;
    wire RU_n_U6052_6;
    wire RXOR0;
    wire RXOR0_n;
    wire RZG_n;
    wand RZ_n;
    wire RZ_n_U5005_4;
    wire RZ_n_U5018_4;
    wire RZ_n_U5051_4;
    wire RZ_n_U6052_2;
    wire S01;
    wire S01_n;
    wire S02;
    wire S02_n;
    wire S03;
    wire S03_n;
    wire S04;
    wire S04_n;
    wire S05;
    wire S05_n;
    wire S06;
    wire S06_n;
    wire S07;
    wire S07_n;
    wire S08;
    wire S08_n;
    wire S09;
    wire S09_n;
    wire S10;
    wire S10_n;
    wire S11;
    wire S11_n;
    wire S12;
    wire S12_n;
    wor SA01;
    wire SA01_U31001_31;
    wire SA01_U31023_16;
    wire SA01_U31025_8;
    wor SA02;
    wire SA02_U31001_33;
    wire SA02_U31023_14;
    wire SA02_U31025_9;
    wor SA03;
    wire SA03_U31001_35;
    wire SA03_U31023_12;
    wire SA03_U31025_10;
    wor SA04;
    wire SA04_U31001_38;
    wire SA04_U31023_9;
    wire SA04_U31025_13;
    wor SA05;
    wire SA05_U31001_40;
    wire SA05_U31023_7;
    wire SA05_U31025_14;
    wor SA06;
    wire SA06_U31001_42;
    wire SA06_U31023_5;
    wire SA06_U31025_15;
    wor SA07;
    wire SA07_U31001_44;
    wire SA07_U31023_3;
    wire SA07_U31025_16;
    wor SA08;
    wire SA08_U31001_30;
    wire SA08_U31024_18;
    wire SA08_U31025_29;
    wor SA09;
    wire SA09_U31001_32;
    wire SA09_U31024_16;
    wire SA09_U31025_30;
    wor SA10;
    wire SA10_U31001_34;
    wire SA10_U31024_14;
    wire SA10_U31025_31;
    wor SA11;
    wire SA11_U31001_36;
    wire SA11_U31024_12;
    wire SA11_U31025_32;
    wor SA12;
    wire SA12_U31001_39;
    wire SA12_U31024_9;
    wire SA12_U31025_35;
    wor SA13;
    wire SA13_U31001_41;
    wire SA13_U31024_7;
    wire SA13_U31025_36;
    wor SA14;
    wire SA14_U31001_43;
    wire SA14_U31024_5;
    wire SA14_U31025_37;
    wor SA16;
    wire SA16_U31001_45;
    wire SA16_U31024_3;
    wire SA16_U31025_38;
    wor SAP;
    wire SAP_U31001_29;
    wire SAP_U31023_18;
    wire SAP_U31025_7;
    wire SB0_n;
    wire SB1_n;
    wire SB2;
    wire SB2_n;
    wire SBE;
    wire SBF;
    wire SBY;
    wand SCAD;
    wire SCAD_U5051_6;
    wire SCAD_U5051_8;
    wire SCAD_n;
    wire SETAB;
    wire SETCD;
    wire SETEK;
    wire SHANC_n;
    wire SHIFT;
    wire SHIFT_n;
    wire SHINC_n;
    wire SQ0_n;
    wire SQ1_n;
    wire SQ2_n;
    wire SQEXT;
    wire SQEXT_n;
    wire SQR10;
    wire SQR10_n;
    wire SQR12_n;
    wire SR_n;
    wire ST0_n;
    wire ST1;
    wire ST1_n;
    wire ST2;
    wand ST2_n;
    wire ST2_n_U5024_6;
    wire ST2_n_U6047_12;
    wire ST3_n;
    wire STBE;
    wire STBF;
    wire STD2;
    wire STFET1_n;
    wire STNDBY_n;
    wire STOP;
    wire STOPA;
    wire STOP_n;
    wire STORE1_n;
    wire STR14;
    wire STR19;
    wire STR210;
    wire STR311;
    wire STR412;
    wire STR58;
    wire STR912;
    wire STRGAT;
    wire STRT1;
    wire STRTFC;
    wire SU0;
    wire SUMA01_n;
    wire SUMA02_n;
    wire SUMA03_n;
    wire SUMA11_n;
    wire SUMA12_n;
    wire SUMA13_n;
    wire SUMA14_n;
    wire SUMA15_n;
    wire SUMA16_n;
    wire SUMB01_n;
    wire SUMB02_n;
    wire SUMB03_n;
    wire SUMB11_n;
    wire SUMB12_n;
    wire SUMB13_n;
    wire SUMB14_n;
    wire SUMB15_n;
    wire SUMB16_n;
    wire T01;
    wire T01_n;
    wire T02;
    wire T02_n;
    wire T03;
    wire T03_n;
    wire T04;
    wire T04_n;
    wire T05;
    wire T05_n;
    wire T06;
    wire T06_n;
    wire T07;
    wire T07_n;
    wire T08;
    wire T08_n;
    wire T09;
    wire T09_n;
    wire T10;
    wire T10_n;
    wire T11;
    wire T11_n;
    wire T12;
    wire T12A;
    wire T12USE_n;
    wire T12_n;
    wire T1P;
    wire T2P;
    wire T3P;
    wire T4P;
    wire T5P;
    wire T6P;
    wire TC0;
    wire TC0_n;
    wire TCF0;
    wire TCSAJ3;
    wire TCSAJ3_n;
    wire THRSTD;
    wire TIMR;
    wire TL15;
    wire TMPOUT;
    wand TMZ_n;
    wire TMZ_n_U4045_12;
    wire TMZ_n_U5012_2;
    wire TMZ_n_U5067_6;
    wand TOV_n;
    wire TOV_n_U5061_2;
    wire TOV_n_U6019_4;
    wire TPARG_n;
    wire TPOR_n;
    wire TPZG_n;
    wire TRSM;
    wire TS0;
    wire TS0_n;
    wand TSGN_n;
    wire TSGN_n_U4063_2;
    wire TSGN_n_U4063_4;
    wire TSGN_n_U5061_12;
    wire TSGN_n_U5067_10;
    wire TSGU_n;
    wire TSUDO_n;
    wire TT_n;
    wire TWOX;
    wire U2BBK;
    wire U2BBKG_n;
    wire UNF_n;
    wire US2SG;
    wire WAG_n;
    wire WALSG_n;
    wire WAND0;
    wand WA_n;
    wire WA_n_U5005_10;
    wire WA_n_U5024_12;
    wire WA_n_U5058_6;
    wire WA_n_U6029_8;
    wire WA_n_U6047_4;
    wire WBBEG_n;
    wire WBG_n;
    wand WB_n;
    wire WB_n_U5018_12;
    wire WB_n_U5041_2;
    wire WB_n_U5041_4;
    wire WB_n_U5061_8;
    wire WB_n_U6014_10;
    wire WCH11_n;
    wire WCHG_n;
    wire WCH_n;
    wire WEBG_n;
    wire WEDOPG_n;
    wire WEX;
    wire WEY;
    wire WFBG_n;
    wire WG1G_n;
    wire WG2G_n;
    wire WG3G_n;
    wire WG4G_n;
    wire WG5G_n;
    wand WG_n;
    wire WG_n_U4039_12;
    wire WG_n_U4045_10;
    wire WG_n_U4045_2;
    wire WG_n_U5012_4;
    wire WG_n_U6019_8;
    wire WG_n_U6037_6;
    wire WHOMP;
    wire WHOMPA;
    wire WL01_n;
    wire WL02_n;
    wire WL03_n;
    wire WL04_n;
    wire WL05_n;
    wire WL06_n;
    wire WL07_n;
    wire WL08_n;
    wire WL09_n;
    wire WL10_n;
    wire WL11_n;
    wire WL12_n;
    wire WL13_n;
    wire WL14_n;
    wire WL15;
    wire WL15_n;
    wire WL16;
    wire WL16_n;
    wire WLG_n;
    wand WL_n;
    wire WL_n_U4061_6;
    wire WL_n_U5067_4;
    wire WL_n_U6014_6;
    wire WOR0;
    wire WOVR_n;
    wire WQG_n;
    wire WQ_n;
    wand WSC_n;
    wire WSC_n_U6019_6;
    wire WSC_n_U6037_4;
    wire WSG_n;
    wand WS_n;
    wire WS_n_U5035_12;
    wire WS_n_U6041_8;
    wire WT;
    wire WT_n;
    wand WY12_n;
    wire WY12_n_U5018_6;
    wire WY12_n_U5046_12;
    wire WYDG_n;
    wire WYDLOG_n;
    wand WYD_n;
    wire WYD_n_U5067_8;
    wire WYD_n_U6004_10;
    wire WYHIG_n;
    wire WYLOG_n;
    wand WY_n;
    wire WY_n_U4061_2;
    wire WY_n_U4061_4;
    wire WY_n_U5012_12;
    wire WY_n_U5024_8;
    wire WY_n_U5046_6;
    wire WY_n_U6004_12;
    wire WZG_n;
    wand WZ_n;
    wire WZ_n_U5018_8;
    wire WZ_n_U5058_12;
    wire WZ_n_U6019_2;
    wire XB0;
    wire XB0_n;
    wire XB1;
    wire XB1E;
    wire XB1_n;
    wire XB2;
    wire XB2E;
    wire XB2_n;
    wire XB3;
    wire XB3E;
    wire XB3_n;
    wire XB4;
    wire XB4E;
    wire XB4_n;
    wire XB5;
    wire XB5E;
    wire XB5_n;
    wire XB6;
    wire XB6E;
    wire XB6_n;
    wire XB7;
    wire XB7E;
    wire XB7_n;
    wire XT0_n;
    wire XT1E;
    wire XT1_n;
    wire XT2E;
    wire XT2_n;
    wire XT3E;
    wire XT3_n;
    wire XT4E;
    wire XT4_n;
    wire XT5E;
    wire XT5_n;
    wire XT6E;
    wire XT6_n;
    wire XT7E;
    wire XUY01_n;
    wire XUY02_n;
    wire XUY05_n;
    wire XUY06_n;
    wire XUY09_n;
    wire XUY10_n;
    wire XUY13_n;
    wire XUY14_n;
    wire YB0_n;
    wire YB1E;
    wire YB2E;
    wire YB3E;
    wire YT0_n;
    wire YT1E;
    wire YT2E;
    wire YT3E;
    wire YT4E;
    wire YT5E;
    wire YT6E;
    wire YT7E;
    wand Z15_n;
    wire Z15_n_U11041_8;
    wire Z15_n_U5067_2;
    wand Z16_n;
    wire Z16_n_U11063_4;
    wire Z16_n_U5058_4;
    wire ZAP_n;
    wire ZID;
    wire ZOUT_n;
    wire __A01_1__CHAT01;
    wire __A01_1__CHAT02;
    wire __A01_1__CHAT03;
    wire __A01_1__CHAT04;
    wire __A01_1__CHAT05;
    wire __A01_1__CHAT06;
    wire __A01_1__CHAT07;
    wire __A01_1__CHAT08;
    wire __A01_1__CHAT09;
    wire __A01_1__CHAT10;
    wire __A01_1__CHAT11;
    wire __A01_1__CHAT12;
    wire __A01_1__F02A;
    wire __A01_1__F02B;
    wire __A01_1__F03A;
    wire __A01_1__F03B;
    wire __A01_1__F05A;
    wire __A01_1__F05B;
    wire __A01_1__F06A;
    wire __A01_1__F08A;
    wire __A01_1__F11A;
    wire __A01_1__F11B;
    wire __A01_1__F12A;
    wire __A01_1__F13A;
    wire __A01_1__F13B;
    wire __A01_1__F14A;
    wire __A01_1__F15A;
    wire __A01_1__F15B;
    wire __A01_1__F16A;
    wire __A01_1__F16B;
    wire __A01_1__FS02;
    wire __A01_1__FS02A;
    wire __A01_1__FS03;
    wire __A01_1__FS03A;
    wire __A01_1__FS04;
    wire __A01_1__FS04A;
    wire __A01_1__FS05;
    wire __A01_1__FS05A;
    wire __A01_1__FS06;
    wire __A01_1__FS07;
    wire __A01_1__FS08;
    wire __A01_1__FS11;
    wire __A01_1__FS12;
    wire __A01_1__FS15;
    wire __A01_1__FS16;
    wire __A01_1__FS17;
    wire __A01_1__scaler_s10__FS_n;
    wire __A01_1__scaler_s11__FS_n;
    wire __A01_1__scaler_s12__FS_n;
    wire __A01_1__scaler_s13__FS_n;
    wire __A01_1__scaler_s14__FS_n;
    wire __A01_1__scaler_s15__FS_n;
    wire __A01_1__scaler_s16__FS_n;
    wire __A01_1__scaler_s17__FS_n;
    wire __A01_1__scaler_s2__FS_n;
    wire __A01_1__scaler_s3__FS_n;
    wire __A01_1__scaler_s4__FS_n;
    wire __A01_1__scaler_s5__FS_n;
    wire __A01_1__scaler_s6__FS_n;
    wire __A01_1__scaler_s7__FS_n;
    wire __A01_1__scaler_s8__FS_n;
    wire __A01_1__scaler_s9__FS_n;
    wire __A01_2__CHAT13;
    wire __A01_2__CHAT14;
    wire __A01_2__CHBT01;
    wire __A01_2__CHBT02;
    wire __A01_2__CHBT03;
    wire __A01_2__CHBT04;
    wire __A01_2__CHBT05;
    wire __A01_2__CHBT06;
    wire __A01_2__CHBT07;
    wire __A01_2__CHBT08;
    wire __A01_2__CHBT09;
    wire __A01_2__CHBT10;
    wire __A01_2__CHBT11;
    wire __A01_2__CHBT12;
    wire __A01_2__CHBT13;
    wire __A01_2__CHBT14;
    wire __A01_2__F18A;
    wire __A01_2__F18B;
    wire __A01_2__F19A;
    wire __A01_2__F19B;
    wire __A01_2__F20A;
    wire __A01_2__F20B;
    wire __A01_2__F21A;
    wire __A01_2__F21B;
    wire __A01_2__F22A;
    wire __A01_2__F22B;
    wire __A01_2__F23A;
    wire __A01_2__F23B;
    wire __A01_2__F24A;
    wire __A01_2__F24B;
    wire __A01_2__F25A;
    wire __A01_2__F25B;
    wire __A01_2__F26A;
    wire __A01_2__F26B;
    wire __A01_2__F27A;
    wire __A01_2__F27B;
    wire __A01_2__F28A;
    wire __A01_2__F28B;
    wire __A01_2__F29A;
    wire __A01_2__F29B;
    wire __A01_2__F30A;
    wire __A01_2__F30B;
    wire __A01_2__F31A;
    wire __A01_2__F31B;
    wire __A01_2__F32A;
    wire __A01_2__F32B;
    wire __A01_2__F33A;
    wire __A01_2__F33B;
    wire __A01_2__FS18;
    wire __A01_2__FS19;
    wire __A01_2__FS20;
    wire __A01_2__FS21;
    wire __A01_2__FS22;
    wire __A01_2__FS23;
    wire __A01_2__FS24;
    wire __A01_2__FS25;
    wire __A01_2__FS26;
    wire __A01_2__FS27;
    wire __A01_2__FS28;
    wire __A01_2__FS29;
    wire __A01_2__FS30;
    wire __A01_2__FS31;
    wire __A01_2__FS32;
    wire __A01_2__FS33;
    wire __A01_2__scaler_s18__FS_n;
    wire __A01_2__scaler_s19__FS_n;
    wire __A01_2__scaler_s20__FS_n;
    wire __A01_2__scaler_s21__FS_n;
    wire __A01_2__scaler_s22__FS_n;
    wire __A01_2__scaler_s23__FS_n;
    wire __A01_2__scaler_s24__FS_n;
    wire __A01_2__scaler_s25__FS_n;
    wire __A01_2__scaler_s26__FS_n;
    wire __A01_2__scaler_s27__FS_n;
    wire __A01_2__scaler_s28__FS_n;
    wire __A01_2__scaler_s29__FS_n;
    wire __A01_2__scaler_s30__FS_n;
    wire __A01_2__scaler_s31__FS_n;
    wire __A01_2__scaler_s32__FS_n;
    wire __A01_2__scaler_s33__FS_n;
    wire __A01_NET_143;
    wire __A01_NET_163;
    wire __A01_NET_177;
    wire __A01_NET_178;
    wire __A01_NET_179;
    wire __A01_NET_180;
    wire __A01_NET_181;
    wire __A01_NET_182;
    wire __A01_NET_183;
    wire __A01_NET_184;
    wire __A01_NET_185;
    wire __A01_NET_186;
    wire __A01_NET_187;
    wire __A01_NET_188;
    wire __A01_NET_189;
    wire __A01_NET_190;
    wire __A01_NET_191;
    wire __A01_NET_192;
    wire __A01_NET_193;
    wire __A01_NET_194;
    wire __A01_NET_195;
    wire __A01_NET_196;
    wire __A01_NET_197;
    wire __A01_NET_198;
    wire __A01_NET_199;
    wire __A01_NET_200;
    wire __A01_NET_201;
    wire __A01_NET_202;
    wire __A01_NET_203;
    wire __A01_NET_204;
    wire __A01_NET_205;
    wire __A01_NET_206;
    wire __A01_NET_207;
    wire __A01_NET_208;
    wire __A01_NET_209;
    wire __A01_NET_210;
    wire __A01_NET_211;
    wire __A01_NET_212;
    wire __A01_NET_213;
    wire __A01_NET_214;
    wire __A01_NET_215;
    wire __A01_NET_216;
    wire __A01_NET_217;
    wire __A01_NET_218;
    wire __A01_NET_219;
    wire __A01_NET_220;
    wire __A01_NET_221;
    wire __A01_NET_222;
    wire __A01_NET_223;
    wire __A01_NET_224;
    wire __A01_NET_225;
    wire __A01_NET_226;
    wire __A01_NET_227;
    wire __A01_NET_228;
    wire __A01_NET_229;
    wire __A01_NET_230;
    wire __A01_NET_231;
    wire __A01_NET_232;
    wire __A01_NET_233;
    wire __A01_NET_234;
    wire __A01_NET_235;
    wire __A01_NET_236;
    wire __A01_NET_237;
    wire __A01_NET_238;
    wire __A01_NET_239;
    wire __A01_NET_240;
    wire __A02_1__EVNSET_n;
    wire __A02_1__ODDSET_n;
    wire __A02_1__OVFSTB_n;
    wire __A02_1__RINGA_n;
    wire __A02_1__RINGB_n;
    wire __A02_1__cdiv_1__A;
    wire __A02_1__cdiv_1__B;
    wire __A02_1__cdiv_1__D;
    wire __A02_1__cdiv_1__FS;
    wire __A02_1__cdiv_1__FS_n;
    wire __A02_1__cdiv_2__A;
    wire __A02_1__cdiv_2__B;
    wire __A02_1__cdiv_2__C;
    wire __A02_1__cdiv_2__D;
    wire __A02_1__cdiv_2__F;
    wire __A02_1__cdiv_2__FS;
    wire __A02_1__cdiv_2__FS_n;
    wire __A02_1__evnset;
    wire __A02_1__oddset;
    wire __A02_1__ovfstb_r1;
    wire __A02_1__ovfstb_r2;
    wire __A02_1__ovfstb_r3;
    wire __A02_1__ovfstb_r4;
    wire __A02_1__ovfstb_r5;
    wire __A02_1__ovfstb_r6;
    wire __A02_2__EDSET;
    wire __A02_2__F01A;
    wire __A02_2__F01B;
    wire __A02_2__F01C;
    wire __A02_2__F01D;
    wire __A02_2__SB0;
    wire __A02_2__SB1;
    wire __A02_2__SB4;
    wire __A02_2__T12DC_n;
    wire __A02_3__OVF;
    wire __A02_3__T01DC_n;
    wire __A02_3__T02DC_n;
    wire __A02_3__T03DC_n;
    wire __A02_3__T04DC_n;
    wire __A02_3__T05DC_n;
    wire __A02_3__T06DC_n;
    wire __A02_3__T07DC_n;
    wire __A02_3__T08DC_n;
    wire __A02_3__T09DC_n;
    wire __A02_3__T10DC_n;
    wand __A02_3__T12SET;
    wire __A02_3__T12SET_U2039_2;
    wire __A02_3__T12SET_U2039_4;
    wire __A02_3__T12SET_U2039_6;
    wire __A02_3__T12SET_U2039_8;
    wire __A02_3__UNF;
    wire __A02_NET_127;
    wire __A02_NET_141;
    wire __A02_NET_142;
    wire __A02_NET_143;
    wire __A02_NET_144;
    wire __A02_NET_145;
    wire __A02_NET_146;
    wire __A02_NET_147;
    wire __A02_NET_148;
    wire __A02_NET_149;
    wire __A02_NET_150;
    wire __A02_NET_151;
    wand __A02_NET_152;
    wire __A02_NET_152_U2020_2;
    wire __A02_NET_152_U2020_4;
    wire __A02_NET_153;
    wire __A02_NET_154;
    wire __A02_NET_155;
    wire __A02_NET_158;
    wire __A02_NET_159;
    wire __A02_NET_160;
    wire __A02_NET_161;
    wire __A02_NET_162;
    wire __A02_NET_163;
    wire __A02_NET_164;
    wire __A02_NET_165;
    wire __A02_NET_166;
    wire __A02_NET_167;
    wire __A02_NET_168;
    wire __A02_NET_169;
    wire __A02_NET_170;
    wire __A02_NET_171;
    wire __A02_NET_172;
    wire __A02_NET_173;
    wire __A02_NET_174;
    wire __A02_NET_175;
    wire __A02_NET_176;
    wire __A02_NET_177;
    wire __A02_NET_178;
    wire __A02_NET_179;
    wire __A02_NET_180;
    wire __A02_NET_181;
    wire __A02_NET_182;
    wire __A02_NET_183;
    wire __A02_NET_184;
    wire __A02_NET_185;
    wire __A02_NET_186;
    wire __A02_NET_187;
    wire __A02_NET_188;
    wire __A02_NET_189;
    wire __A02_NET_190;
    wire __A02_NET_191;
    wire __A02_NET_192;
    wire __A02_NET_193;
    wire __A02_NET_194;
    wire __A02_NET_195;
    wire __A02_NET_196;
    wire __A02_NET_197;
    wire __A02_NET_198;
    wire __A03_1__CSQG;
    wire __A03_1__INHINT;
    wire __A03_1__INKBT1;
    wire __A03_1__MIIP;
    wire __A03_1__MINHL;
    wire __A03_1__MSQ10;
    wire __A03_1__MSQ11;
    wire __A03_1__MSQ12;
    wire __A03_1__MSQ13;
    wire __A03_1__MSQ14;
    wire __A03_1__MSQ16;
    wire __A03_1__MSQEXT;
    wire __A03_1__NISQL;
    wire __A03_1__QC0;
    wire __A03_1__RPTFRC;
    wire __A03_1__SQ3_n;
    wire __A03_1__SQ4_n;
    wire __A03_1__SQ5_n;
    wire __A03_1__SQ6_n;
    wire __A03_1__SQ7_n;
    wire __A03_1__SQR11;
    wire __A03_1__SQR12;
    wire __A03_1__SQR13;
    wire __A03_1__SQR14;
    wire __A03_1__SQR16;
    wire __A03_1__WSQG_n;
    wire __A03_1__wsqg;
    wire __A03_2__AUG0;
    wire __A03_2__BMF0;
    wire __A03_2__BMF0_n;
    wire __A03_2__BZF0;
    wire __A03_2__BZF0_n;
    wire __A03_2__DIM0;
    wand __A03_2__IC13_n;
    wire __A03_2__IC13_n_U3033_2;
    wire __A03_2__IC13_n_U3033_4;
    wire __A03_2__IC3_n;
    wire __A03_2__IC4_n;
    wire __A03_2__IC9_n;
    wire __A03_2__LXCH0;
    wire __A03_2__NDX0;
    wire __A03_2__NDXX1;
    wire __A03_2__NEXST0;
    wire __A03_2__NEXST0_n;
    wire __A03_2__QXCH0;
    wire __A03_2__SQ5QC0_n;
    wire __A03_NET_161;
    wire __A03_NET_163;
    wire __A03_NET_164;
    wire __A03_NET_165;
    wire __A03_NET_166;
    wire __A03_NET_167;
    wire __A03_NET_168;
    wire __A03_NET_169;
    wire __A03_NET_170;
    wire __A03_NET_171;
    wire __A03_NET_172;
    wire __A03_NET_174;
    wire __A03_NET_175;
    wire __A03_NET_176;
    wire __A03_NET_177;
    wire __A03_NET_178;
    wire __A03_NET_179;
    wire __A03_NET_180;
    wire __A03_NET_181;
    wire __A03_NET_182;
    wire __A03_NET_183;
    wire __A03_NET_184;
    wire __A03_NET_185;
    wire __A03_NET_186;
    wire __A03_NET_187;
    wire __A03_NET_188;
    wire __A03_NET_189;
    wire __A03_NET_190;
    wire __A03_NET_191;
    wire __A03_NET_192;
    wire __A03_NET_193;
    wire __A03_NET_194;
    wire __A03_NET_195;
    wire __A03_NET_196;
    wire __A03_NET_197;
    wire __A03_NET_198;
    wire __A03_NET_199;
    wire __A03_NET_200;
    wire __A03_NET_201;
    wire __A03_NET_202;
    wire __A03_NET_203;
    wire __A03_NET_204;
    wire __A03_NET_205;
    wire __A03_NET_206;
    wire __A03_NET_207;
    wire __A03_NET_208;
    wire __A03_NET_209;
    wire __A03_NET_210;
    wire __A03_NET_212;
    wire __A03_NET_213;
    wire __A03_NET_214;
    wire __A03_NET_215;
    wire __A03_NET_216;
    wire __A03_NET_217;
    wire __A03_NET_218;
    wire __A03_NET_219;
    wire __A03_NET_220;
    wire __A03_NET_221;
    wire __A03_NET_225;
    wire __A03_NET_226;
    wire __A03_NET_227;
    wire __A03_NET_229;
    wire __A03_NET_232;
    wire __A03_NET_233;
    wire __A04_1__DV0;
    wire __A04_1__DV0_n;
    wire __A04_1__DV376;
    wire __A04_1__MBR1;
    wire __A04_1__MBR2;
    wire __A04_1__MST1;
    wire __A04_1__MST2;
    wire __A04_1__MST3;
    wand __A04_1__SGUM;
    wire __A04_1__SGUM_U4003_10;
    wire __A04_1__SGUM_U4003_12;
    wire __A04_1__ST1376_n;
    wire __A04_1__ST376;
    wire __A04_1__ST376_n;
    wire __A04_1__ST4_n;
    wire __A04_1__STG1;
    wire __A04_1__STG2;
    wire __A04_1__STG3;
    wire __A04_1__TSGN2;
    wire __A04_2__BR12B;
    wire __A04_2__BR1B2;
    wire __A04_2__BRXP3;
    wire __A04_2__MRSC;
    wire __A04_2__READ0_n;
    wire __A04_2__RUPT0_n;
    wire __A04_2__RUPT1_n;
    wire __A04_2__WOR0_n;
    wire __A04_2__WRITE0;
    wire __A04_2__WRITE0_n;
    wire __A04_NET_185;
    wire __A04_NET_186;
    wire __A04_NET_187;
    wire __A04_NET_188;
    wire __A04_NET_189;
    wire __A04_NET_190;
    wire __A04_NET_191;
    wire __A04_NET_192;
    wire __A04_NET_193;
    wire __A04_NET_194;
    wire __A04_NET_195;
    wire __A04_NET_196;
    wire __A04_NET_197;
    wire __A04_NET_198;
    wire __A04_NET_199;
    wire __A04_NET_200;
    wire __A04_NET_201;
    wire __A04_NET_202;
    wire __A04_NET_203;
    wire __A04_NET_204;
    wire __A04_NET_205;
    wire __A04_NET_208;
    wire __A04_NET_209;
    wire __A04_NET_210;
    wire __A04_NET_211;
    wand __A04_NET_212;
    wire __A04_NET_212_U4029_10;
    wire __A04_NET_212_U4029_8;
    wire __A04_NET_213;
    wand __A04_NET_216;
    wire __A04_NET_216_U4023_2;
    wire __A04_NET_216_U4023_4;
    wand __A04_NET_217;
    wire __A04_NET_217_U4023_6;
    wire __A04_NET_217_U4023_8;
    wire __A04_NET_218;
    wire __A04_NET_219;
    wire __A04_NET_220;
    wire __A04_NET_221;
    wand __A04_NET_222;
    wire __A04_NET_222_U4023_10;
    wire __A04_NET_222_U4023_12;
    wire __A04_NET_222_U4029_2;
    wire __A04_NET_222_U4029_4;
    wire __A04_NET_222_U4029_6;
    wire __A04_NET_229;
    wire __A04_NET_230;
    wire __A04_NET_231;
    wire __A04_NET_232;
    wire __A04_NET_233;
    wire __A04_NET_234;
    wire __A04_NET_235;
    wire __A04_NET_236;
    wire __A04_NET_237;
    wand __A04_NET_238;
    wire __A04_NET_238_U4003_6;
    wire __A04_NET_238_U4003_8;
    wire __A04_NET_241;
    wire __A04_NET_242;
    wire __A04_NET_243;
    wire __A04_NET_244;
    wire __A04_NET_245;
    wire __A04_NET_246;
    wire __A04_NET_247;
    wire __A04_NET_248;
    wire __A04_NET_249;
    wand __A04_NET_250;
    wire __A04_NET_250_U4003_2;
    wire __A04_NET_250_U4003_4;
    wire __A04_NET_251;
    wire __A04_NET_252;
    wire __A04_NET_253;
    wire __A04_NET_254;
    wire __A04_NET_255;
    wire __A04_NET_256;
    wire __A04_NET_259;
    wire __A04_NET_260;
    wire __A04_NET_261;
    wire __A04_NET_262;
    wire __A04_NET_264;
    wire __A04_NET_265;
    wire __A04_NET_266;
    wire __A04_NET_268;
    wire __A04_NET_269;
    wire __A04_NET_270;
    wire __A04_NET_271;
    wire __A04_NET_272;
    wire __A04_NET_273;
    wire __A04_NET_274;
    wire __A04_NET_275;
    wire __A04_NET_276;
    wire __A04_NET_277;
    wire __A04_NET_278;
    wire __A04_NET_279;
    wire __A04_NET_280;
    wire __A04_NET_281;
    wire __A04_NET_282;
    wand __A04_NET_283;
    wire __A04_NET_283_U4045_4;
    wire __A04_NET_283_U4045_6;
    wire __A04_NET_284;
    wire __A04_NET_285;
    wire __A04_NET_286;
    wire __A04_NET_287;
    wire __A04_NET_288;
    wire __A04_NET_289;
    wire __A04_NET_290;
    wire __A04_NET_291;
    wire __A04_NET_292;
    wire __A04_NET_293;
    wire __A04_NET_294;
    wire __A04_NET_295;
    wire __A04_NET_296;
    wire __A04_NET_297;
    wire __A04_NET_298;
    wire __A04_NET_299;
    wire __A04_NET_300;
    wire __A04_NET_302;
    wire __A04_NET_303;
    wire __A04_NET_308;
    wire __A04_NET_309;
    wire __A04_NET_310;
    wire __A04_NET_311;
    wire __A04_NET_312;
    wire __A04_NET_313;
    wire __A04_NET_314;
    wire __A04_NET_315;
    wire __A04_NET_316;
    wire __A04_NET_317;
    wire __A04_NET_318;
    wire __A04_NET_319;
    wire __A04_NET_320;
    wire __A04_NET_321;
    wire __A04_NET_322;
    wire __A04_NET_323;
    wire __A04_NET_324;
    wire __A04_NET_325;
    wire __A04_NET_326;
    wire __A04_NET_327;
    wire __A04_NET_328;
    wire __A04_NET_329;
    wire __A04_NET_330;
    wire __A04_NET_331;
    wire __A04_NET_332;
    wire __A04_NET_335;
    wire __A04_NET_336;
    wire __A04_NET_337;
    wire __A05_1__10XP6;
    wire __A05_1__10XP7;
    wire __A05_1__3XP5;
    wire __A05_1__8XP12;
    wire __A05_1__8XP15;
    wire __A05_1__8XP3;
    wire __A05_1__DV1B1B;
    wire __A05_1__MNISQ;
    wire __A05_1__NISQ_n;
    wire __A05_1__PARTC;
    wire __A05_2__10XP10;
    wire __A05_2__11XP6;
    wire __A05_2__5XP13;
    wire __A05_2__5XP19;
    wire __A05_2__5XP9;
    wire __A05_2__6XP2;
    wire __A05_2__6XP7;
    wire __A05_NET_177;
    wire __A05_NET_178;
    wire __A05_NET_179;
    wire __A05_NET_180;
    wire __A05_NET_181;
    wire __A05_NET_182;
    wire __A05_NET_184;
    wire __A05_NET_185;
    wire __A05_NET_186;
    wire __A05_NET_187;
    wire __A05_NET_188;
    wire __A05_NET_190;
    wire __A05_NET_191;
    wire __A05_NET_193;
    wire __A05_NET_194;
    wire __A05_NET_195;
    wire __A05_NET_196;
    wire __A05_NET_197;
    wire __A05_NET_198;
    wire __A05_NET_199;
    wire __A05_NET_200;
    wire __A05_NET_202;
    wire __A05_NET_203;
    wire __A05_NET_205;
    wire __A05_NET_206;
    wire __A05_NET_207;
    wire __A05_NET_208;
    wire __A05_NET_209;
    wire __A05_NET_212;
    wire __A05_NET_213;
    wire __A05_NET_214;
    wire __A05_NET_215;
    wire __A05_NET_216;
    wire __A05_NET_217;
    wire __A05_NET_218;
    wire __A05_NET_219;
    wire __A05_NET_220;
    wire __A05_NET_221;
    wire __A05_NET_222;
    wire __A05_NET_223;
    wire __A05_NET_224;
    wire __A05_NET_225;
    wire __A05_NET_226;
    wire __A05_NET_227;
    wire __A05_NET_228;
    wire __A05_NET_229;
    wire __A05_NET_230;
    wire __A05_NET_231;
    wire __A05_NET_232;
    wire __A05_NET_233;
    wire __A05_NET_234;
    wire __A05_NET_235;
    wire __A05_NET_236;
    wire __A05_NET_237;
    wire __A05_NET_238;
    wire __A05_NET_239;
    wire __A05_NET_242;
    wire __A05_NET_243;
    wire __A05_NET_244;
    wire __A05_NET_245;
    wire __A05_NET_246;
    wire __A05_NET_247;
    wire __A05_NET_248;
    wire __A05_NET_249;
    wire __A05_NET_250;
    wire __A05_NET_251;
    wire __A05_NET_252;
    wire __A05_NET_253;
    wire __A05_NET_254;
    wire __A05_NET_255;
    wire __A05_NET_256;
    wire __A05_NET_257;
    wire __A05_NET_260;
    wire __A05_NET_261;
    wire __A05_NET_262;
    wire __A05_NET_263;
    wire __A05_NET_264;
    wire __A05_NET_265;
    wire __A05_NET_266;
    wire __A05_NET_268;
    wire __A05_NET_270;
    wire __A05_NET_271;
    wire __A05_NET_272;
    wire __A05_NET_273;
    wire __A05_NET_274;
    wire __A05_NET_275;
    wire __A05_NET_276;
    wire __A05_NET_277;
    wand __A05_NET_278;
    wire __A05_NET_278_U5058_10;
    wire __A05_NET_278_U5058_8;
    wire __A05_NET_279;
    wire __A05_NET_281;
    wire __A05_NET_282;
    wire __A05_NET_283;
    wire __A05_NET_284;
    wire __A05_NET_285;
    wand __A05_NET_287;
    wire __A05_NET_287_U5051_12;
    wire __A05_NET_287_U5058_2;
    wire __A05_NET_288;
    wire __A05_NET_289;
    wire __A05_NET_290;
    wire __A05_NET_291;
    wire __A05_NET_292;
    wire __A05_NET_293;
    wire __A05_NET_294;
    wire __A05_NET_295;
    wire __A05_NET_296;
    wire __A05_NET_297;
    wire __A05_NET_298;
    wand __A05_NET_299;
    wire __A05_NET_299_U5035_10;
    wire __A05_NET_299_U5035_8;
    wire __A05_NET_302;
    wand __A05_NET_303;
    wire __A05_NET_303_U5041_6;
    wire __A05_NET_303_U5041_8;
    wire __A05_NET_304;
    wire __A05_NET_306;
    wire __A05_NET_307;
    wire __A05_NET_308;
    wire __A05_NET_309;
    wire __A05_NET_310;
    wire __A05_NET_311;
    wire __A05_NET_313;
    wire __A05_NET_314;
    wire __A05_NET_315;
    wire __A05_NET_316;
    wire __A05_NET_317;
    wire __A05_NET_319;
    wire __A05_NET_320;
    wire __A05_NET_321;
    wire __A05_NET_322;
    wire __A05_NET_323;
    wire __A05_NET_326;
    wire __A05_NET_327;
    wire __A05_NET_328;
    wire __A05_NET_329;
    wire __A05_NET_330;
    wire __A05_NET_331;
    wire __A05_NET_332;
    wire __A05_NET_333;
    wire __A05_NET_334;
    wire __A05_NET_335;
    wire __A05_NET_336;
    wire __A05_NET_337;
    wire __A05_NET_338;
    wire __A05_NET_339;
    wire __A05_NET_340;
    wire __A05_NET_341;
    wire __A05_NET_342;
    wire __A05_NET_343;
    wire __A05_NET_344;
    wire __A05_NET_345;
    wire __A05_NET_346;
    wire __A05_NET_347;
    wire __A05_NET_349;
    wire __A05_NET_350;
    wire __A05_NET_351;
    wire __A06_1__DVXP1;
    wire __A06_1__L02A_n;
    wire __A06_1__L15A_n;
    wire __A06_1__WHOMP_n;
    wire __A06_1__ZAP;
    wire __A06_1__ZIP;
    wire __A06_1__ZIPCI;
    wire __A06_2__10XP15;
    wire __A06_2__10XP9;
    wire __A06_2__6XP10;
    wire __A06_2__6XP12;
    wire __A06_2__7XP10;
    wire __A06_2__7XP11;
    wire __A06_2__7XP15;
    wire __A06_2__7XP7;
    wire __A06_2__8XP4;
    wire __A06_2__MOUT;
    wire __A06_2__POUT;
    wire __A06_2__RDBANK;
    wire __A06_2__ZOUT;
    wire __A06_NET_181;
    wire __A06_NET_182;
    wire __A06_NET_183;
    wire __A06_NET_184;
    wire __A06_NET_185;
    wire __A06_NET_186;
    wire __A06_NET_188;
    wire __A06_NET_189;
    wire __A06_NET_190;
    wire __A06_NET_191;
    wire __A06_NET_192;
    wire __A06_NET_193;
    wire __A06_NET_195;
    wire __A06_NET_198;
    wire __A06_NET_199;
    wire __A06_NET_200;
    wire __A06_NET_201;
    wire __A06_NET_204;
    wire __A06_NET_205;
    wire __A06_NET_206;
    wire __A06_NET_207;
    wire __A06_NET_208;
    wand __A06_NET_209;
    wire __A06_NET_209_U6041_4;
    wire __A06_NET_209_U6041_6;
    wand __A06_NET_210;
    wire __A06_NET_210_U6041_10;
    wire __A06_NET_210_U6041_12;
    wire __A06_NET_212;
    wire __A06_NET_213;
    wire __A06_NET_214;
    wire __A06_NET_215;
    wire __A06_NET_216;
    wire __A06_NET_217;
    wire __A06_NET_218;
    wire __A06_NET_219;
    wire __A06_NET_221;
    wire __A06_NET_222;
    wire __A06_NET_223;
    wand __A06_NET_224;
    wire __A06_NET_224_U6029_2;
    wire __A06_NET_224_U6029_4;
    wire __A06_NET_225;
    wire __A06_NET_226;
    wire __A06_NET_227;
    wire __A06_NET_228;
    wire __A06_NET_229;
    wire __A06_NET_230;
    wire __A06_NET_231;
    wire __A06_NET_235;
    wire __A06_NET_237;
    wire __A06_NET_238;
    wire __A06_NET_239;
    wire __A06_NET_241;
    wire __A06_NET_243;
    wire __A06_NET_244;
    wire __A06_NET_245;
    wire __A06_NET_246;
    wire __A06_NET_247;
    wand __A06_NET_248;
    wire __A06_NET_248_U6047_10;
    wire __A06_NET_248_U6047_8;
    wire __A06_NET_249;
    wire __A06_NET_250;
    wire __A06_NET_255;
    wire __A06_NET_256;
    wire __A06_NET_257;
    wire __A06_NET_258;
    wire __A06_NET_259;
    wire __A06_NET_262;
    wire __A06_NET_263;
    wire __A06_NET_264;
    wire __A06_NET_265;
    wire __A06_NET_266;
    wire __A06_NET_267;
    wand __A06_NET_268;
    wire __A06_NET_268_U6019_10;
    wire __A06_NET_268_U6019_12;
    wire __A06_NET_269;
    wire __A06_NET_270;
    wire __A06_NET_271;
    wire __A06_NET_272;
    wire __A06_NET_274;
    wire __A06_NET_276;
    wire __A06_NET_277;
    wire __A06_NET_278;
    wire __A06_NET_279;
    wire __A06_NET_280;
    wire __A06_NET_281;
    wire __A06_NET_282;
    wire __A06_NET_283;
    wand __A06_NET_284;
    wire __A06_NET_284_U6014_2;
    wire __A06_NET_284_U6014_4;
    wire __A06_NET_285;
    wire __A06_NET_286;
    wire __A06_NET_287;
    wire __A06_NET_288;
    wire __A06_NET_289;
    wire __A06_NET_290;
    wand __A06_NET_291;
    wire __A06_NET_291_U6004_2;
    wire __A06_NET_291_U6004_4;
    wire __A06_NET_292;
    wire __A06_NET_293;
    wire __A06_NET_294;
    wire __A06_NET_295;
    wire __A06_NET_296;
    wire __A06_NET_301;
    wire __A06_NET_302;
    wire __A06_NET_303;
    wire __A06_NET_304;
    wire __A06_NET_305;
    wire __A06_NET_306;
    wire __A06_NET_307;
    wire __A06_NET_308;
    wire __A06_NET_309;
    wire __A06_NET_310;
    wire __A06_NET_311;
    wire __A06_NET_313;
    wire __A06_NET_314;
    wire __A06_NET_315;
    wire __A06_NET_316;
    wire __A06_NET_317;
    wire __A06_NET_318;
    wire __A06_NET_319;
    wire __A06_NET_320;
    wire __A06_NET_321;
    wire __A06_NET_322;
    wire __A06_NET_323;
    wire __A06_NET_324;
    wire __A06_NET_325;
    wire __A06_NET_326;
    wire __A06_NET_327;
    wire __A06_NET_328;
    wire __A06_NET_329;
    wire __A06_NET_330;
    wire __A06_NET_331;
    wire __A06_NET_332;
    wire __A06_NET_333;
    wire __A06_NET_334;
    wire __A06_NET_335;
    wire __A06_NET_340;
    wire __A06_NET_342;
    wire __A06_NET_343;
    wire __A06_NET_344;
    wire __A06_NET_345;
    wire __A06_NET_346;
    wire __A06_NET_347;
    wire __A06_NET_348;
    wire __A06_NET_349;
    wire __A06_NET_350;
    wire __A07_1__MWAG;
    wire __A07_1__MWBG;
    wire __A07_1__MWG;
    wire __A07_1__MWLG;
    wire __A07_1__MWQG;
    wire __A07_1__MWSG;
    wire __A07_1__MWYG;
    wire __A07_1__MWZG;
    wire __A07_1__P04A;
    wire __A07_1__PIPSAM_n;
    wire __A07_1__WALSG;
    wire __A07_1__WGA_n;
    wire __A07_1__WGNORM;
    wire __A07_1__WSCG_n;
    wire __A07_2__CIFF;
    wire __A07_2__CINORM;
    wire __A07_2__G2LSG;
    wire __A07_2__MRAG;
    wire __A07_2__MRGG;
    wire __A07_2__MRLG;
    wire __A07_2__MRULOG;
    wire __A07_2__MWBBEG;
    wire __A07_2__MWEBG;
    wire __A07_2__MWFBG;
    wire __A07_2__RBBK;
    wire __A07_2__RCHG_n;
    wire __A07_2__RSCG_n;
    wire __A07_2__RUSG_n;
    wire __A07_NET_137;
    wire __A07_NET_138;
    wire __A07_NET_139;
    wire __A07_NET_140;
    wire __A07_NET_141;
    wire __A07_NET_142;
    wire __A07_NET_145;
    wire __A07_NET_148;
    wire __A07_NET_149;
    wire __A07_NET_151;
    wire __A07_NET_152;
    wire __A07_NET_153;
    wire __A07_NET_154;
    wire __A07_NET_155;
    wire __A07_NET_156;
    wire __A07_NET_157;
    wire __A07_NET_158;
    wire __A07_NET_159;
    wire __A07_NET_160;
    wire __A07_NET_161;
    wand __A07_NET_162;
    wire __A07_NET_162_U7007_2;
    wire __A07_NET_162_U7007_4;
    wire __A07_NET_163;
    wire __A07_NET_164;
    wire __A07_NET_165;
    wire __A07_NET_166;
    wire __A07_NET_167;
    wire __A07_NET_168;
    wire __A07_NET_169;
    wire __A07_NET_170;
    wire __A07_NET_171;
    wire __A07_NET_172;
    wire __A07_NET_173;
    wire __A07_NET_174;
    wire __A07_NET_175;
    wire __A07_NET_177;
    wire __A07_NET_178;
    wire __A07_NET_179;
    wire __A07_NET_180;
    wire __A07_NET_181;
    wire __A07_NET_182;
    wire __A07_NET_183;
    wire __A07_NET_184;
    wire __A07_NET_185;
    wire __A07_NET_186;
    wire __A07_NET_187;
    wire __A07_NET_188;
    wire __A07_NET_189;
    wire __A07_NET_190;
    wire __A07_NET_191;
    wire __A07_NET_192;
    wire __A07_NET_194;
    wire __A07_NET_195;
    wire __A07_NET_198;
    wire __A07_NET_199;
    wire __A07_NET_201;
    wire __A07_NET_202;
    wire __A07_NET_203;
    wire __A07_NET_204;
    wire __A07_NET_205;
    wire __A07_NET_206;
    wire __A07_NET_207;
    wire __A07_NET_208;
    wire __A07_NET_209;
    wire __A07_NET_210;
    wire __A07_NET_211;
    wire __A07_NET_212;
    wire __A07_NET_213;
    wire __A07_NET_215;
    wire __A08_1__X1;
    wire __A08_1__X1_n;
    wire __A08_1__X2;
    wire __A08_1__X2_n;
    wire __A08_1__Y1;
    wire __A08_1__Y1_n;
    wire __A08_1__Y2;
    wire __A08_1__Y2_n;
    wire __A08_1___A1_n;
    wire __A08_1___A2_n;
    wire __A08_1___B1_n;
    wire __A08_1___B2_n;
    wire __A08_1___CI_INTERNAL;
    wand __A08_1___G2_n;
    wire __A08_1___G2_n_U8028_10;
    wire __A08_1___G2_n_U8028_12;
    wire __A08_1___MWL1;
    wire __A08_1___MWL2;
    wire __A08_1___Q1_n;
    wire __A08_1___Q2_n;
    wire __A08_1___RL_OUT_1;
    wire __A08_1___RL_OUT_2;
    wire __A08_1___WL1;
    wire __A08_1___WL2;
    wand __A08_1___Z1_n;
    wire __A08_1___Z1_n_U8007_8;
    wand __A08_1___Z2_n;
    wire __A08_1___Z2_n_U8028_4;
    wire __A08_2__X1;
    wire __A08_2__X1_n;
    wire __A08_2__X2;
    wire __A08_2__X2_n;
    wire __A08_2__Y1;
    wire __A08_2__Y1_n;
    wire __A08_2__Y2;
    wire __A08_2__Y2_n;
    wire __A08_2___A1_n;
    wire __A08_2___A2_n;
    wire __A08_2___B1_n;
    wire __A08_2___B2_n;
    wire __A08_2___CI_IN;
    wire __A08_2___CI_INTERNAL;
    wand __A08_2___CO_IN;
    wire __A08_2___CO_IN_U8007_2;
    wire __A08_2___CO_IN_U8013_2;
    wand __A08_2___G1_n;
    wire __A08_2___G1_n_U8050_6;
    wire __A08_2___G1_n_U8050_8;
    wand __A08_2___G2_n;
    wire __A08_2___G2_n_U8063_10;
    wire __A08_2___G2_n_U8063_12;
    wand __A08_2___L1_n;
    wire __A08_2___L1_n_U8041_6;
    wire __A08_2___MWL1;
    wire __A08_2___MWL2;
    wire __A08_2___Q1_n;
    wire __A08_2___Q2_n;
    wire __A08_2___RL_OUT_1;
    wire __A08_2___RL_OUT_2;
    wire __A08_2___SUMA2;
    wire __A08_2___SUMB2;
    wire __A08_2___WL1;
    wire __A08_2___WL2;
    wire __A08_2___XUY1;
    wire __A08_2___XUY2;
    wand __A08_2___Z1_n;
    wire __A08_2___Z1_n_U8041_8;
    wand __A08_2___Z2_n;
    wire __A08_2___Z2_n_U8063_4;
    wire __A08_NET_137;
    wire __A08_NET_138;
    wire __A08_NET_139;
    wire __A08_NET_140;
    wire __A08_NET_141;
    wire __A08_NET_142;
    wire __A08_NET_143;
    wire __A08_NET_144;
    wire __A08_NET_145;
    wire __A08_NET_146;
    wire __A08_NET_147;
    wire __A08_NET_148;
    wire __A08_NET_149;
    wire __A08_NET_152;
    wire __A08_NET_155;
    wire __A08_NET_156;
    wire __A08_NET_157;
    wire __A08_NET_158;
    wire __A08_NET_159;
    wire __A08_NET_160;
    wire __A08_NET_161;
    wire __A08_NET_162;
    wire __A08_NET_163;
    wire __A08_NET_164;
    wire __A08_NET_167;
    wire __A08_NET_168;
    wire __A08_NET_169;
    wire __A08_NET_170;
    wire __A08_NET_175;
    wire __A08_NET_176;
    wire __A08_NET_177;
    wire __A08_NET_178;
    wire __A08_NET_179;
    wire __A08_NET_180;
    wire __A08_NET_181;
    wire __A08_NET_182;
    wire __A08_NET_183;
    wire __A08_NET_184;
    wire __A08_NET_185;
    wire __A08_NET_186;
    wire __A08_NET_187;
    wire __A08_NET_188;
    wire __A08_NET_189;
    wire __A08_NET_190;
    wire __A08_NET_191;
    wire __A08_NET_192;
    wire __A08_NET_193;
    wire __A08_NET_194;
    wire __A08_NET_195;
    wire __A08_NET_196;
    wire __A08_NET_197;
    wire __A08_NET_198;
    wire __A08_NET_199;
    wire __A08_NET_200;
    wire __A08_NET_205;
    wire __A08_NET_206;
    wire __A08_NET_207;
    wire __A08_NET_209;
    wire __A08_NET_210;
    wire __A08_NET_211;
    wire __A08_NET_212;
    wire __A08_NET_213;
    wire __A08_NET_214;
    wire __A08_NET_215;
    wire __A08_NET_216;
    wire __A08_NET_219;
    wire __A08_NET_220;
    wire __A08_NET_221;
    wire __A08_NET_222;
    wire __A08_NET_223;
    wire __A08_NET_224;
    wire __A08_NET_225;
    wire __A08_NET_226;
    wire __A08_NET_227;
    wire __A08_NET_228;
    wire __A08_NET_229;
    wire __A08_NET_230;
    wire __A08_NET_231;
    wire __A08_NET_232;
    wire __A08_NET_233;
    wire __A08_NET_234;
    wire __A08_NET_235;
    wire __A08_NET_236;
    wire __A08_NET_237;
    wire __A08_NET_238;
    wire __A08_NET_239;
    wire __A08_NET_240;
    wire __A08_NET_241;
    wire __A08_NET_242;
    wire __A08_NET_245;
    wire __A08_NET_248;
    wire __A08_NET_249;
    wire __A08_NET_250;
    wire __A08_NET_251;
    wire __A08_NET_252;
    wire __A08_NET_253;
    wire __A08_NET_254;
    wire __A08_NET_255;
    wire __A08_NET_256;
    wire __A08_NET_257;
    wire __A08_NET_260;
    wire __A08_NET_261;
    wire __A08_NET_262;
    wire __A08_NET_263;
    wire __A08_NET_268;
    wire __A08_NET_269;
    wire __A08_NET_270;
    wire __A08_NET_271;
    wire __A08_NET_272;
    wire __A08_NET_273;
    wire __A08_NET_274;
    wire __A08_NET_275;
    wire __A08_NET_276;
    wire __A08_NET_277;
    wire __A08_NET_278;
    wire __A08_NET_279;
    wire __A08_NET_280;
    wire __A08_NET_281;
    wire __A08_NET_282;
    wire __A08_NET_283;
    wire __A08_NET_284;
    wire __A08_NET_285;
    wire __A08_NET_286;
    wire __A08_NET_287;
    wire __A08_NET_288;
    wire __A08_NET_289;
    wire __A08_NET_290;
    wire __A08_NET_291;
    wire __A08_NET_293;
    wire __A08_NET_294;
    wire __A08_NET_298;
    wire __A08_NET_299;
    wire __A08_NET_300;
    wire __A08_NET_302;
    wire __A08_NET_303;
    wire __A08_NET_304;
    wire __A08_NET_305;
    wire __A08_NET_306;
    wire __A08_NET_307;
    wire __A08_NET_308;
    wire __A08_NET_309;
    wire __A08_NET_312;
    wire __A08_NET_313;
    wire __A08_NET_314;
    wire __A08_NET_315;
    wire __A08_NET_316;
    wire __A08_NET_317;
    wire __A08_NET_318;
    wire __A08_NET_319;
    wire __A08_NET_320;
    wire __A08_NET_321;
    wire __A08_NET_322;
    wire __A09_1__X1;
    wire __A09_1__X1_n;
    wire __A09_1__X2;
    wire __A09_1__X2_n;
    wire __A09_1__Y1;
    wire __A09_1__Y1_n;
    wire __A09_1__Y2;
    wire __A09_1__Y2_n;
    wire __A09_1___A1_n;
    wire __A09_1___A2_n;
    wire __A09_1___B1_n;
    wire __A09_1___B2_n;
    wire __A09_1___CI_INTERNAL;
    wand __A09_1___L1_n;
    wire __A09_1___L1_n_U9007_6;
    wand __A09_1___L2_n;
    wire __A09_1___L2_n_U9013_12;
    wire __A09_1___MWL1;
    wire __A09_1___MWL2;
    wire __A09_1___Q1_n;
    wire __A09_1___Q2_n;
    wire __A09_1___RL_OUT_1;
    wire __A09_1___RL_OUT_2;
    wire __A09_1___SUMA1;
    wire __A09_1___SUMA2;
    wire __A09_1___SUMB1;
    wire __A09_1___SUMB2;
    wire __A09_1___WL1;
    wire __A09_1___WL2;
    wand __A09_1___Z1_n;
    wire __A09_1___Z1_n_U9007_8;
    wand __A09_1___Z2_n;
    wire __A09_1___Z2_n_U9028_4;
    wire __A09_2__X1;
    wire __A09_2__X1_n;
    wire __A09_2__X2;
    wire __A09_2__X2_n;
    wire __A09_2__Y1;
    wire __A09_2__Y1_n;
    wire __A09_2__Y2;
    wire __A09_2__Y2_n;
    wire __A09_2___A1_n;
    wire __A09_2___A2_n;
    wire __A09_2___B1_n;
    wire __A09_2___B2_n;
    wire __A09_2___CI_IN;
    wire __A09_2___CI_INTERNAL;
    wand __A09_2___CO_IN;
    wire __A09_2___CO_IN_U9007_2;
    wire __A09_2___CO_IN_U9013_2;
    wand __A09_2___G2_n;
    wire __A09_2___G2_n_U9063_10;
    wire __A09_2___G2_n_U9063_12;
    wand __A09_2___L1_n;
    wire __A09_2___L1_n_U9041_6;
    wire __A09_2___MWL1;
    wire __A09_2___MWL2;
    wire __A09_2___Q1_n;
    wire __A09_2___Q2_n;
    wand __A09_2___RL1_n;
    wire __A09_2___RL1_n_U9041_10;
    wire __A09_2___RL1_n_U9041_12;
    wire __A09_2___RL1_n_U9041_4;
    wire __A09_2___RL1_n_U9050_4;
    wand __A09_2___RL2_n;
    wire __A09_2___RL2_n_U9050_10;
    wire __A09_2___RL2_n_U9063_2;
    wire __A09_2___RL2_n_U9063_6;
    wire __A09_2___RL2_n_U9063_8;
    wire __A09_2___RL_OUT_1;
    wire __A09_2___RL_OUT_2;
    wire __A09_2___SUMA1;
    wire __A09_2___SUMA2;
    wire __A09_2___SUMB1;
    wire __A09_2___SUMB2;
    wire __A09_2___WL1;
    wire __A09_2___WL2;
    wire __A09_2___XUY1;
    wire __A09_2___XUY2;
    wand __A09_2___Z1_n;
    wire __A09_2___Z1_n_U9041_8;
    wand __A09_2___Z2_n;
    wire __A09_2___Z2_n_U9063_4;
    wire __A09_NET_130;
    wire __A09_NET_131;
    wire __A09_NET_132;
    wire __A09_NET_133;
    wire __A09_NET_134;
    wire __A09_NET_135;
    wire __A09_NET_136;
    wire __A09_NET_137;
    wire __A09_NET_138;
    wire __A09_NET_139;
    wire __A09_NET_140;
    wire __A09_NET_141;
    wire __A09_NET_142;
    wire __A09_NET_145;
    wire __A09_NET_148;
    wire __A09_NET_149;
    wire __A09_NET_150;
    wire __A09_NET_151;
    wire __A09_NET_152;
    wire __A09_NET_153;
    wire __A09_NET_154;
    wire __A09_NET_155;
    wire __A09_NET_156;
    wire __A09_NET_157;
    wire __A09_NET_160;
    wire __A09_NET_161;
    wire __A09_NET_162;
    wire __A09_NET_163;
    wire __A09_NET_168;
    wire __A09_NET_169;
    wire __A09_NET_170;
    wire __A09_NET_171;
    wire __A09_NET_172;
    wire __A09_NET_173;
    wire __A09_NET_174;
    wire __A09_NET_175;
    wire __A09_NET_176;
    wire __A09_NET_177;
    wire __A09_NET_178;
    wire __A09_NET_179;
    wire __A09_NET_180;
    wire __A09_NET_181;
    wire __A09_NET_182;
    wire __A09_NET_183;
    wire __A09_NET_184;
    wire __A09_NET_185;
    wire __A09_NET_186;
    wire __A09_NET_187;
    wire __A09_NET_188;
    wire __A09_NET_189;
    wire __A09_NET_190;
    wire __A09_NET_191;
    wire __A09_NET_192;
    wire __A09_NET_193;
    wire __A09_NET_198;
    wire __A09_NET_199;
    wire __A09_NET_200;
    wire __A09_NET_202;
    wire __A09_NET_203;
    wire __A09_NET_204;
    wire __A09_NET_205;
    wire __A09_NET_206;
    wire __A09_NET_207;
    wire __A09_NET_208;
    wire __A09_NET_209;
    wire __A09_NET_212;
    wire __A09_NET_213;
    wire __A09_NET_214;
    wire __A09_NET_215;
    wire __A09_NET_216;
    wire __A09_NET_217;
    wire __A09_NET_218;
    wire __A09_NET_219;
    wire __A09_NET_220;
    wire __A09_NET_221;
    wire __A09_NET_222;
    wire __A09_NET_223;
    wire __A09_NET_224;
    wire __A09_NET_225;
    wire __A09_NET_226;
    wire __A09_NET_227;
    wire __A09_NET_228;
    wire __A09_NET_229;
    wire __A09_NET_230;
    wire __A09_NET_231;
    wire __A09_NET_232;
    wire __A09_NET_233;
    wire __A09_NET_234;
    wire __A09_NET_235;
    wire __A09_NET_238;
    wire __A09_NET_241;
    wire __A09_NET_242;
    wire __A09_NET_243;
    wire __A09_NET_244;
    wire __A09_NET_245;
    wire __A09_NET_246;
    wire __A09_NET_247;
    wire __A09_NET_248;
    wire __A09_NET_249;
    wire __A09_NET_250;
    wire __A09_NET_253;
    wire __A09_NET_254;
    wire __A09_NET_255;
    wire __A09_NET_256;
    wire __A09_NET_261;
    wire __A09_NET_262;
    wire __A09_NET_263;
    wire __A09_NET_264;
    wire __A09_NET_265;
    wire __A09_NET_266;
    wire __A09_NET_267;
    wire __A09_NET_268;
    wire __A09_NET_269;
    wire __A09_NET_270;
    wire __A09_NET_271;
    wire __A09_NET_272;
    wire __A09_NET_273;
    wire __A09_NET_274;
    wire __A09_NET_275;
    wire __A09_NET_276;
    wire __A09_NET_277;
    wire __A09_NET_278;
    wire __A09_NET_279;
    wire __A09_NET_280;
    wire __A09_NET_281;
    wire __A09_NET_282;
    wire __A09_NET_283;
    wire __A09_NET_284;
    wire __A09_NET_286;
    wire __A09_NET_287;
    wire __A09_NET_291;
    wire __A09_NET_292;
    wire __A09_NET_293;
    wire __A09_NET_295;
    wire __A09_NET_296;
    wire __A09_NET_297;
    wire __A09_NET_298;
    wire __A09_NET_299;
    wire __A09_NET_300;
    wire __A09_NET_301;
    wire __A09_NET_302;
    wire __A09_NET_305;
    wire __A09_NET_306;
    wire __A09_NET_307;
    wire __A09_NET_308;
    wire __A09_NET_309;
    wire __A09_NET_310;
    wire __A09_NET_311;
    wire __A09_NET_312;
    wire __A09_NET_313;
    wire __A09_NET_314;
    wire __A09_NET_315;
    wire __A10_1__X1;
    wire __A10_1__X1_n;
    wire __A10_1__X2;
    wire __A10_1__X2_n;
    wire __A10_1__Y1;
    wire __A10_1__Y1_n;
    wire __A10_1__Y2;
    wire __A10_1__Y2_n;
    wire __A10_1___A1_n;
    wire __A10_1___A2_n;
    wire __A10_1___B1_n;
    wire __A10_1___B2_n;
    wire __A10_1___CI_INTERNAL;
    wand __A10_1___L1_n;
    wire __A10_1___L1_n_U10007_6;
    wand __A10_1___L2_n;
    wire __A10_1___L2_n_U10013_12;
    wire __A10_1___MWL1;
    wire __A10_1___MWL2;
    wire __A10_1___Q1_n;
    wire __A10_1___Q2_n;
    wire __A10_1___RL_OUT_1;
    wire __A10_1___RL_OUT_2;
    wire __A10_1___SUMA1;
    wire __A10_1___SUMA2;
    wire __A10_1___SUMB1;
    wire __A10_1___SUMB2;
    wire __A10_1___WL1;
    wire __A10_1___WL2;
    wand __A10_1___Z1_n;
    wire __A10_1___Z1_n_U10007_8;
    wand __A10_1___Z2_n;
    wire __A10_1___Z2_n_U10028_4;
    wire __A10_2__X1;
    wire __A10_2__X1_n;
    wire __A10_2__X2;
    wire __A10_2__X2_n;
    wire __A10_2__Y1;
    wire __A10_2__Y1_n;
    wire __A10_2__Y2;
    wire __A10_2__Y2_n;
    wire __A10_2___A1_n;
    wire __A10_2___A2_n;
    wire __A10_2___B1_n;
    wire __A10_2___B2_n;
    wire __A10_2___CI_IN;
    wire __A10_2___CI_INTERNAL;
    wand __A10_2___CO_IN;
    wire __A10_2___CO_IN_U10007_2;
    wire __A10_2___CO_IN_U10013_2;
    wand __A10_2___G2_n;
    wire __A10_2___G2_n_U10063_10;
    wire __A10_2___G2_n_U10063_12;
    wand __A10_2___L1_n;
    wire __A10_2___L1_n_U10041_6;
    wire __A10_2___MWL1;
    wire __A10_2___MWL2;
    wire __A10_2___Q1_n;
    wire __A10_2___Q2_n;
    wire __A10_2___RL_OUT_1;
    wire __A10_2___RL_OUT_2;
    wire __A10_2___WL1;
    wire __A10_2___WL2;
    wire __A10_2___XUY1;
    wire __A10_2___XUY2;
    wand __A10_2___Z1_n;
    wire __A10_2___Z1_n_U10041_8;
    wand __A10_2___Z2_n;
    wire __A10_2___Z2_n_U10063_4;
    wire __A10_NET_129;
    wire __A10_NET_130;
    wire __A10_NET_131;
    wire __A10_NET_132;
    wire __A10_NET_133;
    wire __A10_NET_134;
    wire __A10_NET_135;
    wire __A10_NET_136;
    wire __A10_NET_137;
    wire __A10_NET_138;
    wire __A10_NET_139;
    wire __A10_NET_140;
    wire __A10_NET_141;
    wire __A10_NET_144;
    wire __A10_NET_147;
    wire __A10_NET_148;
    wire __A10_NET_149;
    wire __A10_NET_150;
    wire __A10_NET_151;
    wire __A10_NET_152;
    wire __A10_NET_153;
    wire __A10_NET_154;
    wire __A10_NET_155;
    wire __A10_NET_156;
    wire __A10_NET_159;
    wire __A10_NET_160;
    wire __A10_NET_161;
    wire __A10_NET_162;
    wire __A10_NET_167;
    wire __A10_NET_168;
    wire __A10_NET_169;
    wire __A10_NET_170;
    wire __A10_NET_171;
    wire __A10_NET_172;
    wire __A10_NET_173;
    wire __A10_NET_174;
    wire __A10_NET_175;
    wire __A10_NET_176;
    wire __A10_NET_177;
    wire __A10_NET_178;
    wire __A10_NET_179;
    wire __A10_NET_180;
    wire __A10_NET_181;
    wire __A10_NET_182;
    wire __A10_NET_183;
    wire __A10_NET_184;
    wire __A10_NET_185;
    wire __A10_NET_186;
    wire __A10_NET_187;
    wire __A10_NET_188;
    wire __A10_NET_189;
    wire __A10_NET_190;
    wire __A10_NET_191;
    wire __A10_NET_192;
    wire __A10_NET_197;
    wire __A10_NET_198;
    wire __A10_NET_199;
    wire __A10_NET_201;
    wire __A10_NET_202;
    wire __A10_NET_203;
    wire __A10_NET_204;
    wire __A10_NET_205;
    wire __A10_NET_206;
    wire __A10_NET_207;
    wire __A10_NET_208;
    wire __A10_NET_211;
    wire __A10_NET_212;
    wire __A10_NET_213;
    wire __A10_NET_214;
    wire __A10_NET_215;
    wire __A10_NET_216;
    wire __A10_NET_217;
    wire __A10_NET_218;
    wire __A10_NET_219;
    wire __A10_NET_220;
    wire __A10_NET_221;
    wire __A10_NET_222;
    wire __A10_NET_223;
    wire __A10_NET_224;
    wire __A10_NET_225;
    wire __A10_NET_226;
    wire __A10_NET_227;
    wire __A10_NET_228;
    wire __A10_NET_229;
    wire __A10_NET_230;
    wire __A10_NET_231;
    wire __A10_NET_232;
    wire __A10_NET_233;
    wire __A10_NET_234;
    wire __A10_NET_237;
    wire __A10_NET_240;
    wire __A10_NET_241;
    wire __A10_NET_242;
    wire __A10_NET_243;
    wire __A10_NET_244;
    wire __A10_NET_245;
    wire __A10_NET_246;
    wire __A10_NET_247;
    wire __A10_NET_248;
    wire __A10_NET_249;
    wire __A10_NET_252;
    wire __A10_NET_253;
    wire __A10_NET_254;
    wire __A10_NET_255;
    wire __A10_NET_260;
    wire __A10_NET_261;
    wire __A10_NET_262;
    wire __A10_NET_263;
    wire __A10_NET_264;
    wire __A10_NET_265;
    wire __A10_NET_266;
    wire __A10_NET_267;
    wire __A10_NET_268;
    wire __A10_NET_269;
    wire __A10_NET_270;
    wire __A10_NET_271;
    wire __A10_NET_272;
    wire __A10_NET_273;
    wire __A10_NET_274;
    wire __A10_NET_275;
    wire __A10_NET_276;
    wire __A10_NET_277;
    wire __A10_NET_278;
    wire __A10_NET_279;
    wire __A10_NET_280;
    wire __A10_NET_281;
    wire __A10_NET_282;
    wire __A10_NET_283;
    wire __A10_NET_285;
    wire __A10_NET_286;
    wire __A10_NET_290;
    wire __A10_NET_291;
    wire __A10_NET_292;
    wire __A10_NET_294;
    wire __A10_NET_295;
    wire __A10_NET_296;
    wire __A10_NET_297;
    wire __A10_NET_298;
    wire __A10_NET_299;
    wire __A10_NET_300;
    wire __A10_NET_301;
    wire __A10_NET_304;
    wire __A10_NET_305;
    wire __A10_NET_306;
    wire __A10_NET_307;
    wire __A10_NET_308;
    wire __A10_NET_309;
    wire __A10_NET_310;
    wire __A10_NET_311;
    wire __A10_NET_312;
    wire __A10_NET_313;
    wire __A10_NET_314;
    wire __A11_1__X1;
    wire __A11_1__X1_n;
    wire __A11_1__X2;
    wire __A11_1__X2_n;
    wire __A11_1__Y1;
    wire __A11_1__Y1_n;
    wire __A11_1__Y2;
    wire __A11_1__Y2_n;
    wire __A11_1___A1_n;
    wire __A11_1___A2_n;
    wire __A11_1___B1_n;
    wire __A11_1___B2_n;
    wire __A11_1___CI_INTERNAL;
    wand __A11_1___L1_n;
    wire __A11_1___L1_n_U11007_6;
    wand __A11_1___L2_n;
    wire __A11_1___L2_n_U11013_12;
    wire __A11_1___MWL1;
    wire __A11_1___MWL2;
    wire __A11_1___Q1_n;
    wire __A11_1___Q2_n;
    wire __A11_1___RL_OUT_1;
    wire __A11_1___RL_OUT_2;
    wire __A11_1___WL1;
    wire __A11_1___WL2;
    wand __A11_1___Z1_n;
    wire __A11_1___Z1_n_U11007_8;
    wand __A11_1___Z2_n;
    wire __A11_1___Z2_n_U11028_4;
    wire __A11_2__X1;
    wire __A11_2__X1_n;
    wire __A11_2__X2;
    wire __A11_2__X2_n;
    wire __A11_2__Y1;
    wire __A11_2__Y1_n;
    wire __A11_2__Y2;
    wire __A11_2__Y2_n;
    wire __A11_2___A1_n;
    wire __A11_2___A2_n;
    wire __A11_2___B1_n;
    wire __A11_2___B2_n;
    wire __A11_2___CI_IN;
    wire __A11_2___CI_INTERNAL;
    wand __A11_2___CO_IN;
    wire __A11_2___CO_IN_U11007_2;
    wire __A11_2___CO_IN_U11013_2;
    wand __A11_2___CO_OUT;
    wire __A11_2___CO_OUT_U11041_2;
    wire __A11_2___CO_OUT_U11050_2;
    wand __A11_2___G2_n;
    wire __A11_2___G2_n_U11063_10;
    wire __A11_2___G2_n_U11063_12;
    wire __A11_2___GEM1;
    wire __A11_2___MWL1;
    wire __A11_2___MWL2;
    wire __A11_2___Q1_n;
    wire __A11_2___Q2_n;
    wire __A11_2___RL_OUT_1;
    wire __A11_2___RL_OUT_2;
    wire __A11_2___XUY1;
    wire __A11_2___XUY2;
    wire __A11_NET_130;
    wire __A11_NET_131;
    wire __A11_NET_132;
    wire __A11_NET_133;
    wire __A11_NET_134;
    wire __A11_NET_135;
    wire __A11_NET_136;
    wire __A11_NET_137;
    wire __A11_NET_138;
    wire __A11_NET_139;
    wire __A11_NET_140;
    wire __A11_NET_141;
    wire __A11_NET_142;
    wire __A11_NET_145;
    wire __A11_NET_148;
    wire __A11_NET_149;
    wire __A11_NET_150;
    wire __A11_NET_151;
    wire __A11_NET_152;
    wire __A11_NET_153;
    wire __A11_NET_154;
    wire __A11_NET_155;
    wire __A11_NET_156;
    wire __A11_NET_157;
    wire __A11_NET_160;
    wire __A11_NET_161;
    wire __A11_NET_162;
    wire __A11_NET_163;
    wire __A11_NET_168;
    wire __A11_NET_169;
    wire __A11_NET_170;
    wire __A11_NET_171;
    wire __A11_NET_172;
    wire __A11_NET_173;
    wire __A11_NET_174;
    wire __A11_NET_175;
    wire __A11_NET_176;
    wire __A11_NET_177;
    wire __A11_NET_178;
    wire __A11_NET_179;
    wire __A11_NET_180;
    wire __A11_NET_181;
    wire __A11_NET_182;
    wire __A11_NET_183;
    wire __A11_NET_184;
    wire __A11_NET_185;
    wire __A11_NET_186;
    wire __A11_NET_187;
    wire __A11_NET_188;
    wire __A11_NET_189;
    wire __A11_NET_190;
    wire __A11_NET_191;
    wire __A11_NET_192;
    wire __A11_NET_193;
    wire __A11_NET_198;
    wire __A11_NET_199;
    wire __A11_NET_200;
    wire __A11_NET_202;
    wire __A11_NET_203;
    wire __A11_NET_204;
    wire __A11_NET_205;
    wire __A11_NET_206;
    wire __A11_NET_207;
    wire __A11_NET_208;
    wire __A11_NET_209;
    wire __A11_NET_212;
    wire __A11_NET_213;
    wire __A11_NET_214;
    wire __A11_NET_215;
    wire __A11_NET_216;
    wire __A11_NET_217;
    wire __A11_NET_218;
    wire __A11_NET_219;
    wire __A11_NET_220;
    wire __A11_NET_221;
    wire __A11_NET_222;
    wire __A11_NET_223;
    wire __A11_NET_224;
    wire __A11_NET_225;
    wire __A11_NET_226;
    wire __A11_NET_227;
    wire __A11_NET_228;
    wire __A11_NET_229;
    wire __A11_NET_230;
    wire __A11_NET_231;
    wire __A11_NET_232;
    wire __A11_NET_233;
    wire __A11_NET_234;
    wire __A11_NET_235;
    wire __A11_NET_238;
    wire __A11_NET_241;
    wire __A11_NET_242;
    wire __A11_NET_243;
    wire __A11_NET_244;
    wire __A11_NET_245;
    wire __A11_NET_246;
    wire __A11_NET_247;
    wire __A11_NET_248;
    wire __A11_NET_249;
    wire __A11_NET_250;
    wire __A11_NET_253;
    wire __A11_NET_254;
    wire __A11_NET_255;
    wire __A11_NET_256;
    wire __A11_NET_261;
    wire __A11_NET_262;
    wire __A11_NET_263;
    wire __A11_NET_264;
    wire __A11_NET_265;
    wire __A11_NET_266;
    wire __A11_NET_267;
    wire __A11_NET_268;
    wire __A11_NET_269;
    wire __A11_NET_270;
    wire __A11_NET_271;
    wire __A11_NET_272;
    wire __A11_NET_273;
    wire __A11_NET_274;
    wire __A11_NET_275;
    wire __A11_NET_276;
    wire __A11_NET_277;
    wire __A11_NET_278;
    wire __A11_NET_279;
    wire __A11_NET_280;
    wire __A11_NET_281;
    wire __A11_NET_282;
    wire __A11_NET_283;
    wire __A11_NET_284;
    wire __A11_NET_286;
    wire __A11_NET_287;
    wire __A11_NET_291;
    wire __A11_NET_292;
    wire __A11_NET_293;
    wire __A11_NET_295;
    wire __A11_NET_296;
    wire __A11_NET_297;
    wire __A11_NET_298;
    wire __A11_NET_299;
    wire __A11_NET_300;
    wire __A11_NET_301;
    wire __A11_NET_302;
    wire __A11_NET_305;
    wire __A11_NET_306;
    wire __A11_NET_307;
    wire __A11_NET_308;
    wire __A11_NET_309;
    wire __A11_NET_310;
    wire __A11_NET_311;
    wire __A11_NET_312;
    wire __A11_NET_313;
    wire __A11_NET_314;
    wire __A11_NET_315;
    wire __A12_1__G01A_n;
    wire __A12_1__G02_n;
    wire __A12_1__G03_n;
    wire __A12_1__G16A_n;
    wand __A12_1__GNZRO;
    wire __A12_1__GNZRO_U12016_2;
    wire __A12_1__GNZRO_U12016_4;
    wire __A12_1__MGP_n;
    wire __A12_1__MPAL;
    wire __A12_1__MSP;
    wire __A12_1__PA03;
    wire __A12_1__PA03_n;
    wire __A12_1__PA06;
    wire __A12_1__PA06_n;
    wire __A12_1__PA09;
    wire __A12_1__PA09_n;
    wire __A12_1__PA12;
    wire __A12_1__PA12_n;
    wire __A12_1__PA15;
    wire __A12_1__PA15_n;
    wire __A12_1__PB09;
    wire __A12_1__PB09_n;
    wire __A12_1__PB15;
    wire __A12_1__PB15_n;
    wire __A12_1__PC15;
    wire __A12_1__T7PHS4;
    wire __A12_1__T7PHS4_n;
    wire __A12_2__G01A;
    wire __A12_NET_110;
    wire __A12_NET_113;
    wire __A12_NET_114;
    wire __A12_NET_115;
    wire __A12_NET_116;
    wire __A12_NET_117;
    wire __A12_NET_119;
    wire __A12_NET_121;
    wire __A12_NET_122;
    wire __A12_NET_123;
    wire __A12_NET_124;
    wire __A12_NET_125;
    wire __A12_NET_126;
    wire __A12_NET_127;
    wire __A12_NET_128;
    wire __A12_NET_129;
    wire __A12_NET_130;
    wire __A12_NET_131;
    wire __A12_NET_132;
    wire __A12_NET_133;
    wire __A12_NET_134;
    wire __A12_NET_135;
    wire __A12_NET_136;
    wire __A12_NET_137;
    wire __A12_NET_138;
    wire __A12_NET_139;
    wire __A12_NET_140;
    wire __A12_NET_141;
    wire __A12_NET_142;
    wire __A12_NET_143;
    wire __A12_NET_144;
    wire __A12_NET_145;
    wire __A12_NET_146;
    wire __A12_NET_147;
    wire __A12_NET_150;
    wire __A12_NET_151;
    wire __A12_NET_152;
    wire __A12_NET_153;
    wire __A12_NET_154;
    wire __A12_NET_155;
    wire __A12_NET_158;
    wire __A12_NET_163;
    wire __A12_NET_170;
    wire __A12_NET_171;
    wire __A12_NET_177;
    wire __A12_NET_180;
    wire __A12_NET_181;
    wire __A12_NET_184;
    wire __A12_NET_185;
    wire __A12_NET_186;
    wire __A12_NET_187;
    wire __A12_NET_190;
    wire __A12_NET_191;
    wire __A12_NET_192;
    wire __A12_NET_193;
    wire __A12_NET_194;
    wire __A12_NET_195;
    wire __A12_NET_196;
    wire __A12_NET_197;
    wire __A12_NET_198;
    wire __A12_NET_199;
    wire __A12_NET_200;
    wire __A12_NET_201;
    wire __A12_NET_207;
    wire __A12_NET_208;
    wire __A12_NET_209;
    wire __A12_NET_210;
    wire __A12_NET_211;
    wire __A12_NET_212;
    wire __A12_NET_213;
    wire __A12_NET_214;
    wire __A12_NET_215;
    wire __A12_NET_216;
    wire __A12_NET_217;
    wire __A12_NET_218;
    wire __A12_NET_219;
    wire __A12_NET_220;
    wire __A12_NET_221;
    wire __A12_NET_222;
    wire __A12_NET_223;
    wire __A12_NET_224;
    wire __A12_NET_225;
    wire __A12_NET_226;
    wire __A12_NET_227;
    wire __A12_NET_228;
    wire __A12_NET_229;
    wire __A12_NET_230;
    wire __A12_NET_231;
    wire __A12_NET_232;
    wire __A12_NET_233;
    wire __A12_NET_234;
    wire __A12_NET_235;
    wire __A12_NET_236;
    wire __A12_NET_237;
    wire __A12_NET_238;
    wire __A12_NET_239;
    wire __A12_NET_240;
    wire __A12_NET_241;
    wire __A12_NET_242;
    wire __A12_NET_243;
    wire __A12_NET_244;
    wire __A12_NET_245;
    wire __A12_NET_246;
    wire __A12_NET_248;
    wire __A12_NET_249;
    wire __A12_NET_250;
    wire __A12_NET_251;
    wire __A12_NET_254;
    wire __A12_NET_255;
    wire __A12_NET_256;
    wire __A12_NET_257;
    wire __A13_1__CGCWAR;
    wand __A13_1__CKTAL_n;
    wire __A13_1__CKTAL_n_U13006_2;
    wire __A13_1__CKTAL_n_U13006_4;
    wire __A13_1__CON1;
    wire __A13_1__CON2;
    wire __A13_1__CON3;
    wire __A13_1__DOFILT;
    wire __A13_1__F12B_n;
    wire __A13_1__F14H;
    wire __A13_1__FILTIN;
    wire __A13_1__FS13_n;
    wire __A13_1__MCTRAL_n;
    wire __A13_1__MOSCAL_n;
    wire __A13_1__MPIPAL_n;
    wire __A13_1__MRPTAL_n;
    wire __A13_1__MSCAFL_n;
    wire __A13_1__MSCDBL_n;
    wire __A13_1__MTCAL_n;
    wire __A13_1__MVFAIL_n;
    wire __A13_1__MWARNF_n;
    wire __A13_1__MWATCH_n;
    wire __A13_1__NOTEST;
    wire __A13_1__NOTEST_n;
    wire __A13_1__RESTRT;
    wire __A13_1__SBYEXT;
    wire __A13_1__SCADBL;
    wire __A13_1__SYNC14_n;
    wire __A13_1__SYNC4_n;
    wire __A13_1__TMPCAU;
    wire __A13_1__WARN;
    wire __A13_1__WATCH;
    wire __A13_1__WATCHP;
    wire __A13_2__INOTRD;
    wire __A13_2__MINKL;
    wire __A13_2__MREQIN;
    wire __A13_2__STORE1;
    wire __A13_NET_158;
    wire __A13_NET_159;
    wire __A13_NET_160;
    wire __A13_NET_161;
    wire __A13_NET_162;
    wire __A13_NET_163;
    wire __A13_NET_164;
    wire __A13_NET_166;
    wire __A13_NET_167;
    wire __A13_NET_168;
    wire __A13_NET_169;
    wire __A13_NET_170;
    wire __A13_NET_171;
    wire __A13_NET_175;
    wire __A13_NET_178;
    wire __A13_NET_179;
    wire __A13_NET_180;
    wire __A13_NET_181;
    wand __A13_NET_182;
    wire __A13_NET_182_U13021_2;
    wire __A13_NET_182_U13021_4;
    wire __A13_NET_187;
    wire __A13_NET_188;
    wire __A13_NET_189;
    wire __A13_NET_192;
    wire __A13_NET_193;
    wire __A13_NET_197;
    wire __A13_NET_198;
    wire __A13_NET_199;
    wire __A13_NET_200;
    wire __A13_NET_202;
    wire __A13_NET_206;
    wire __A13_NET_207;
    wire __A13_NET_208;
    wire __A13_NET_209;
    wire __A13_NET_210;
    wire __A13_NET_213;
    wire __A13_NET_214;
    wire __A13_NET_219;
    wire __A13_NET_220;
    wire __A13_NET_221;
    wire __A13_NET_222;
    wire __A13_NET_223;
    wire __A13_NET_226;
    wire __A13_NET_227;
    wire __A13_NET_228;
    wire __A13_NET_229;
    wire __A13_NET_230;
    wire __A13_NET_231;
    wire __A13_NET_232;
    wire __A13_NET_233;
    wire __A13_NET_234;
    wire __A13_NET_235;
    wire __A13_NET_236;
    wire __A13_NET_237;
    wire __A13_NET_238;
    wire __A13_NET_243;
    wire __A13_NET_244;
    wire __A13_NET_249;
    wire __A13_NET_250;
    wire __A13_NET_251;
    wire __A13_NET_252;
    wire __A13_NET_253;
    wire __A13_NET_254;
    wire __A13_NET_255;
    wire __A13_NET_257;
    wire __A13_NET_258;
    wire __A13_NET_259;
    wire __A13_NET_260;
    wire __A13_NET_261;
    wire __A13_NET_262;
    wire __A13_NET_263;
    wire __A13_NET_264;
    wire __A13_NET_265;
    wand __A13_NET_266;
    wire __A13_NET_266_U13006_10;
    wire __A13_NET_266_U13006_12;
    wire __A13_NET_266_U13006_6;
    wire __A13_NET_266_U13006_8;
    wire __A13_NET_266_U13021_10;
    wire __A13_NET_266_U13021_12;
    wire __A13_NET_266_U13021_6;
    wire __A13_NET_266_U13021_8;
    wire __A13_NET_266_U13036_2;
    wire __A13_NET_266_U13036_4;
    wire __A13_NET_266_U13036_6;
    wire __A13_NET_267;
    wire __A13_NET_268;
    wire __A13_NET_270;
    wire __A13_NET_272;
    wire __A13_NET_273;
    wire __A13_NET_274;
    wire __A13_NET_275;
    wire __A13_NET_276;
    wire __A13_NET_277;
    wire __A13_NET_280;
    wire __A13_NET_281;
    wire __A13_NET_284;
    wire __A13_NET_285;
    wire __A13_NET_286;
    wire __A13_NET_287;
    wire __A13_NET_288;
    wire __A13_NET_289;
    wire __A13_NET_290;
    wire __A13_NET_291;
    wire __A13_NET_292;
    wire __A13_NET_293;
    wire __A13_NET_294;
    wire __A13_NET_297;
    wire __A13_NET_298;
    wire __A13_NET_299;
    wire __A13_NET_300;
    wire __A13_NET_301;
    wire __A13_NET_302;
    wand __A13_NET_303;
    wire __A13_NET_303_U13036_10;
    wire __A13_NET_303_U13036_8;
    wire __A13_NET_304;
    wire __A13_NET_305;
    wire __A13_NET_306;
    wire __A13_NET_307;
    wire __A13_NET_308;
    wire __A13_NET_309;
    wire __A13_NET_310;
    wire __A13_NET_311;
    wire __A13_NET_312;
    wire __A13_NET_313;
    wire __A14_1__CLEARA;
    wire __A14_1__CLEARB;
    wire __A14_1__CLEARC;
    wire __A14_1__CLEARD;
    wand __A14_1__ERAS;
    wire __A14_1__ERAS_U14014_10;
    wire __A14_1__ERAS_U14014_12;
    wire __A14_1__ERAS_n;
    wire __A14_1__FNERAS_n;
    wire __A14_1__IHENV;
    wire __A14_1__REDRST;
    wire __A14_1__REX;
    wire __A14_1__REY;
    wire __A14_1__ROP_n;
    wire __A14_1__RSTKX_n;
    wire __A14_1__RSTKY_n;
    wire __A14_1__RSTK_n;
    wire __A14_1__S08A;
    wire __A14_1__S08A_n;
    wire __A14_1__SBESET;
    wand __A14_1__SBFSET;
    wire __A14_1__SBFSET_U14014_2;
    wire __A14_1__SBFSET_U14014_4;
    wire __A14_1__SETAB_n;
    wire __A14_1__SETCD_n;
    wand __A14_1__TPGE;
    wire __A14_1__TPGE_U14033_2;
    wire __A14_1__TPGE_U14033_4;
    wand __A14_1__TPGF;
    wire __A14_1__TPGF_U14014_6;
    wire __A14_1__TPGF_U14014_8;
    wire __A14_2__EAD09;
    wire __A14_2__EAD09_n;
    wire __A14_2__EAD10;
    wire __A14_2__EAD10_n;
    wire __A14_2__EAD11;
    wire __A14_2__EAD11_n;
    wire __A14_2__IL01_n;
    wire __A14_2__IL02_n;
    wire __A14_2__IL03_n;
    wire __A14_2__IL04_n;
    wire __A14_2__IL05_n;
    wire __A14_2__IL06_n;
    wire __A14_2__IL07_n;
    wire __A14_2__ILP;
    wire __A14_2__ILP_n;
    wire __A14_2__RILP1;
    wire __A14_2__RILP1_n;
    wire __A14_2__XB0E;
    wire __A14_2__XT0;
    wire __A14_2__XT0E;
    wire __A14_2__XT1;
    wire __A14_2__XT2;
    wire __A14_2__XT3;
    wire __A14_2__XT4;
    wire __A14_2__XT5;
    wire __A14_2__XT6;
    wire __A14_2__XT7;
    wire __A14_2__XT7_n;
    wire __A14_2__YB0;
    wire __A14_2__YB0E;
    wire __A14_2__YB1;
    wire __A14_2__YB1_n;
    wire __A14_2__YB2;
    wire __A14_2__YB2_n;
    wire __A14_2__YB3;
    wire __A14_2__YB3_n;
    wire __A14_2__YT0;
    wire __A14_2__YT0E;
    wire __A14_2__YT1;
    wire __A14_2__YT1_n;
    wire __A14_2__YT2;
    wire __A14_2__YT2_n;
    wire __A14_2__YT3;
    wire __A14_2__YT3_n;
    wire __A14_2__YT4;
    wire __A14_2__YT4_n;
    wire __A14_2__YT5;
    wire __A14_2__YT5_n;
    wire __A14_2__YT6;
    wire __A14_2__YT6_n;
    wire __A14_2__YT7;
    wire __A14_2__YT7_n;
    wire __A14_NET_192;
    wire __A14_NET_194;
    wire __A14_NET_196;
    wire __A14_NET_198;
    wire __A14_NET_199;
    wire __A14_NET_200;
    wire __A14_NET_202;
    wire __A14_NET_203;
    wire __A14_NET_204;
    wire __A14_NET_205;
    wire __A14_NET_206;
    wire __A14_NET_207;
    wire __A14_NET_208;
    wire __A14_NET_209;
    wire __A14_NET_210;
    wire __A14_NET_211;
    wire __A14_NET_212;
    wire __A14_NET_213;
    wire __A14_NET_214;
    wire __A14_NET_215;
    wire __A14_NET_216;
    wire __A14_NET_217;
    wire __A14_NET_218;
    wire __A14_NET_219;
    wire __A14_NET_220;
    wire __A14_NET_221;
    wire __A14_NET_222;
    wire __A14_NET_223;
    wire __A14_NET_224;
    wire __A14_NET_225;
    wire __A14_NET_226;
    wire __A14_NET_231;
    wire __A14_NET_232;
    wire __A14_NET_233;
    wire __A14_NET_234;
    wire __A14_NET_235;
    wire __A14_NET_236;
    wire __A14_NET_237;
    wire __A14_NET_238;
    wire __A14_NET_239;
    wire __A14_NET_240;
    wire __A14_NET_241;
    wire __A14_NET_242;
    wire __A14_NET_246;
    wire __A14_NET_247;
    wire __A14_NET_248;
    wire __A14_NET_249;
    wire __A14_NET_250;
    wire __A14_NET_251;
    wire __A14_NET_252;
    wire __A14_NET_253;
    wire __A14_NET_254;
    wire __A14_NET_255;
    wire __A14_NET_256;
    wire __A14_NET_257;
    wire __A14_NET_258;
    wire __A14_NET_259;
    wire __A14_NET_260;
    wire __A14_NET_261;
    wire __A14_NET_262;
    wire __A14_NET_263;
    wire __A14_NET_264;
    wire __A14_NET_265;
    wire __A14_NET_266;
    wire __A14_NET_267;
    wire __A14_NET_268;
    wire __A14_NET_269;
    wire __A14_NET_270;
    wire __A14_NET_271;
    wire __A14_NET_272;
    wire __A14_NET_274;
    wire __A14_NET_275;
    wire __A14_NET_276;
    wire __A14_NET_279;
    wire __A14_NET_280;
    wire __A14_NET_285;
    wire __A14_NET_286;
    wire __A14_NET_287;
    wire __A14_NET_288;
    wire __A14_NET_289;
    wire __A14_NET_290;
    wire __A14_NET_292;
    wire __A14_NET_295;
    wire __A14_NET_296;
    wire __A14_NET_297;
    wire __A14_NET_300;
    wire __A14_NET_301;
    wire __A14_NET_306;
    wire __A14_NET_308;
    wire __A15_1__BBK1;
    wire __A15_1__BBK2;
    wire __A15_1__BBK3;
    wire __A15_1__BK16;
    wire __A15_1__DNRPTA;
    wire __A15_1__EB10_n;
    wire __A15_1__EB11;
    wire __A15_1__EB9_n;
    wire __A15_1__F11;
    wire __A15_1__F11_n;
    wire __A15_1__F12;
    wire __A15_1__F12_n;
    wire __A15_1__F13;
    wire __A15_1__F13_n;
    wire __A15_1__F14;
    wire __A15_1__F14_n;
    wire __A15_1__F15;
    wire __A15_1__F15_n;
    wire __A15_1__F16;
    wire __A15_1__F16_n;
    wire __A15_1__FB11;
    wire __A15_1__FB11_n;
    wire __A15_1__FB12;
    wire __A15_1__FB12_n;
    wire __A15_1__FB13;
    wire __A15_1__FB13_n;
    wire __A15_1__FB14;
    wire __A15_1__FB14_n;
    wire __A15_1__FB16;
    wire __A15_1__FB16_n;
    wire __A15_1__KRPTA_n;
    wire __A15_1__PRPOR1;
    wire __A15_1__PRPOR2;
    wire __A15_1__PRPOR3;
    wire __A15_1__PRPOR4;
    wire __A15_1__RPTA12;
    wire __A15_1__RPTAD6;
    wire __A15_1__RRPA1_n;
    wire __A15_2__036H;
    wire __A15_2__036L;
    wire __A15_2__147H;
    wire __A15_2__147L;
    wire __A15_2__2510H;
    wire __A15_2__2510L;
    wire __A15_2__KY1RST;
    wire __A15_2__KY2RST;
    wire __A15_2__NE00;
    wire __A15_2__NE01;
    wire __A15_2__NE012_n;
    wire __A15_2__NE02;
    wire __A15_2__NE03;
    wire __A15_2__NE036_n;
    wire __A15_2__NE04;
    wire __A15_2__NE05;
    wire __A15_2__NE06;
    wire __A15_2__NE07;
    wire __A15_2__NE10;
    wire __A15_2__NE147_n;
    wire __A15_2__NE2510_n;
    wire __A15_2__NE345_n;
    wire __A15_2__NE6710_n;
    wire __A15_2__RPTAD3;
    wire __A15_2__RPTAD4;
    wire __A15_2__RPTAD5;
    wire __A15_2__T6RPT;
    wire __A15_NET_149;
    wire __A15_NET_150;
    wire __A15_NET_151;
    wire __A15_NET_152;
    wire __A15_NET_153;
    wire __A15_NET_154;
    wire __A15_NET_155;
    wire __A15_NET_156;
    wire __A15_NET_157;
    wire __A15_NET_158;
    wire __A15_NET_159;
    wire __A15_NET_160;
    wire __A15_NET_161;
    wire __A15_NET_162;
    wire __A15_NET_163;
    wire __A15_NET_164;
    wire __A15_NET_165;
    wire __A15_NET_166;
    wire __A15_NET_167;
    wire __A15_NET_168;
    wire __A15_NET_169;
    wire __A15_NET_170;
    wire __A15_NET_171;
    wire __A15_NET_172;
    wire __A15_NET_173;
    wire __A15_NET_174;
    wire __A15_NET_175;
    wire __A15_NET_176;
    wire __A15_NET_179;
    wire __A15_NET_180;
    wire __A15_NET_183;
    wire __A15_NET_184;
    wire __A15_NET_185;
    wire __A15_NET_189;
    wire __A15_NET_191;
    wire __A15_NET_192;
    wire __A15_NET_193;
    wire __A15_NET_194;
    wire __A15_NET_195;
    wire __A15_NET_196;
    wire __A15_NET_197;
    wire __A15_NET_198;
    wire __A15_NET_199;
    wire __A15_NET_200;
    wire __A15_NET_202;
    wire __A15_NET_203;
    wire __A15_NET_204;
    wire __A15_NET_205;
    wire __A15_NET_212;
    wire __A15_NET_213;
    wire __A15_NET_214;
    wire __A15_NET_215;
    wire __A15_NET_216;
    wire __A15_NET_217;
    wire __A15_NET_218;
    wire __A15_NET_219;
    wire __A15_NET_220;
    wire __A15_NET_221;
    wire __A15_NET_222;
    wire __A15_NET_223;
    wire __A15_NET_224;
    wire __A15_NET_225;
    wire __A15_NET_226;
    wire __A15_NET_227;
    wire __A15_NET_228;
    wire __A15_NET_229;
    wand __A15_NET_230;
    wire __A15_NET_230_U15016_12;
    wire __A15_NET_230_U15039_2;
    wire __A15_NET_231;
    wire __A15_NET_232;
    wire __A15_NET_233;
    wire __A15_NET_234;
    wire __A15_NET_235;
    wire __A15_NET_236;
    wand __A15_NET_237;
    wire __A15_NET_237_U15016_10;
    wire __A15_NET_237_U15016_8;
    wire __A15_NET_245;
    wire __A15_NET_246;
    wire __A15_NET_252;
    wire __A15_NET_253;
    wire __A15_NET_254;
    wire __A15_NET_255;
    wire __A15_NET_256;
    wire __A15_NET_257;
    wire __A15_NET_258;
    wire __A15_NET_260;
    wire __A15_NET_261;
    wire __A15_NET_263;
    wire __A15_NET_270;
    wire __A15_NET_273;
    wire __A15_NET_274;
    wire __A15_NET_276;
    wire __A15_NET_277;
    wire __A15_NET_278;
    wire __A15_NET_279;
    wire __A15_NET_280;
    wire __A15_NET_281;
    wire __A15_NET_282;
    wire __A15_NET_284;
    wire __A15_NET_285;
    wire __A15_NET_286;
    wire __A15_NET_287;
    wire __A15_NET_288;
    wire __A15_NET_289;
    wire __A15_NET_290;
    wire __A15_NET_291;
    wire __A15_NET_292;
    wire __A15_NET_293;
    wire __A15_NET_294;
    wire __A15_NET_295;
    wire __A15_NET_296;
    wire __A15_NET_298;
    wire __A15_NET_301;
    wire __A15_NET_302;
    wire __A15_NET_304;
    wire __A15_NET_305;
    wire __A15_NET_306;
    wire __A15_NET_307;
    wire __A15_NET_308;
    wire __A16_1__CCH05;
    wire __A16_1__CCH06;
    wire __A16_1__CCH12;
    wire __A16_1__CH1207;
    wire __A16_1__CH1208;
    wand __A16_1__CHOR01_n;
    wire __A16_1__CHOR01_n_U16004_2;
    wand __A16_1__CHOR02_n;
    wire __A16_1__CHOR02_n_U16004_4;
    wand __A16_1__CHOR03_n;
    wire __A16_1__CHOR03_n_U16004_6;
    wand __A16_1__CHOR04_n;
    wire __A16_1__CHOR04_n_U16004_8;
    wand __A16_1__CHOR05_n;
    wire __A16_1__CHOR05_n_U16004_10;
    wand __A16_1__CHOR06_n;
    wire __A16_1__CHOR06_n_U16004_12;
    wand __A16_1__CHOR07_n;
    wire __A16_1__CHOR07_n_U16021_2;
    wand __A16_1__CHOR08_n;
    wire __A16_1__CHOR08_n_U16021_4;
    wire __A16_1__OT1207;
    wire __A16_1__OT1207_n;
    wire __A16_1__RCH05_n;
    wire __A16_1__RCH06_n;
    wire __A16_1__RCH12_n;
    wire __A16_1__RCmXmP;
    wire __A16_1__RCmXmY;
    wire __A16_1__RCmXpP;
    wire __A16_1__RCmXpY;
    wire __A16_1__RCmYmR;
    wire __A16_1__RCmYpR;
    wire __A16_1__RCmZmR;
    wire __A16_1__RCmZpR;
    wire __A16_1__RCpXmP;
    wire __A16_1__RCpXmY;
    wire __A16_1__RCpXpP;
    wire __A16_1__RCpXpY;
    wire __A16_1__RCpYmR;
    wire __A16_1__RCpYpR;
    wire __A16_1__RCpZmR;
    wire __A16_1__RCpZpR;
    wire __A16_1__TVCNAB;
    wire __A16_1__WCH05_n;
    wire __A16_1__WCH06_n;
    wire __A16_1__WCH12_n;
    wire __A16_2__CH1209;
    wire __A16_2__CH1210;
    wire __A16_2__CH1211;
    wire __A16_2__CH1212;
    wand __A16_2__CHOR01_n;
    wire __A16_2__CHOR01_n_U16021_6;
    wand __A16_2__CHOR02_n;
    wire __A16_2__CHOR02_n_U16021_8;
    wand __A16_2__CHOR03_n;
    wire __A16_2__CHOR03_n_U16021_10;
    wand __A16_2__CHOR04_n;
    wire __A16_2__CHOR04_n_U16021_12;
    wand __A16_2__CHOR05_n;
    wire __A16_2__CHOR05_n_U16044_2;
    wand __A16_2__CHOR06_n;
    wire __A16_2__CHOR06_n_U16044_4;
    wand __A16_2__CHOR07_n;
    wire __A16_2__CHOR07_n_U16044_6;
    wire __A16_2__COARSE;
    wire __A16_2__COMACT;
    wire __A16_2__DISDAC;
    wire __A16_2__ENERIM;
    wire __A16_2__ENEROP;
    wire __A16_2__KYRLS;
    wire __A16_2__MROLGT;
    wire __A16_2__OPEROR;
    wire __A16_2__S4BOFF;
    wire __A16_2__S4BSEQ;
    wire __A16_2__S4BTAK;
    wire __A16_2__STARON;
    wire __A16_2__UPLACT;
    wire __A16_2__VNFLSH;
    wire __A16_2__ZEROPT;
    wire __A16_2__ZIMCDU;
    wire __A16_2__ZOPCDU;
    wire __A16_NET_108;
    wire __A16_NET_109;
    wire __A16_NET_110;
    wire __A16_NET_111;
    wire __A16_NET_112;
    wire __A16_NET_113;
    wire __A16_NET_114;
    wire __A16_NET_115;
    wire __A16_NET_116;
    wire __A16_NET_117;
    wire __A16_NET_118;
    wire __A16_NET_119;
    wire __A16_NET_120;
    wire __A16_NET_121;
    wire __A16_NET_122;
    wire __A16_NET_123;
    wire __A16_NET_124;
    wire __A16_NET_125;
    wire __A16_NET_126;
    wire __A16_NET_127;
    wire __A16_NET_128;
    wire __A16_NET_129;
    wire __A16_NET_130;
    wire __A16_NET_131;
    wire __A16_NET_132;
    wire __A16_NET_133;
    wire __A16_NET_134;
    wire __A16_NET_135;
    wire __A16_NET_136;
    wire __A16_NET_137;
    wire __A16_NET_138;
    wire __A16_NET_139;
    wire __A16_NET_140;
    wire __A16_NET_141;
    wire __A16_NET_142;
    wire __A16_NET_143;
    wire __A16_NET_144;
    wire __A16_NET_145;
    wire __A16_NET_146;
    wire __A16_NET_147;
    wire __A16_NET_148;
    wire __A16_NET_149;
    wire __A16_NET_150;
    wire __A16_NET_151;
    wire __A16_NET_152;
    wire __A16_NET_153;
    wire __A16_NET_154;
    wire __A16_NET_155;
    wire __A16_NET_156;
    wire __A16_NET_157;
    wire __A16_NET_158;
    wire __A16_NET_159;
    wire __A16_NET_160;
    wire __A16_NET_161;
    wire __A16_NET_162;
    wire __A16_NET_163;
    wire __A16_NET_167;
    wire __A16_NET_168;
    wire __A16_NET_169;
    wire __A16_NET_170;
    wire __A16_NET_171;
    wire __A16_NET_172;
    wire __A16_NET_174;
    wire __A16_NET_177;
    wire __A16_NET_178;
    wire __A16_NET_179;
    wire __A16_NET_180;
    wire __A16_NET_181;
    wire __A16_NET_182;
    wire __A16_NET_183;
    wire __A16_NET_184;
    wire __A16_NET_185;
    wire __A16_NET_186;
    wire __A16_NET_187;
    wire __A16_NET_188;
    wire __A16_NET_189;
    wire __A16_NET_190;
    wire __A16_NET_191;
    wire __A16_NET_192;
    wire __A16_NET_193;
    wire __A16_NET_194;
    wire __A16_NET_195;
    wire __A16_NET_196;
    wire __A16_NET_197;
    wire __A16_NET_198;
    wire __A16_NET_199;
    wire __A16_NET_200;
    wire __A16_NET_201;
    wire __A16_NET_202;
    wire __A16_NET_203;
    wire __A16_NET_204;
    wire __A16_NET_205;
    wire __A16_NET_206;
    wire __A16_NET_207;
    wire __A16_NET_208;
    wire __A16_NET_209;
    wire __A16_NET_210;
    wire __A16_NET_211;
    wire __A16_NET_212;
    wire __A16_NET_213;
    wire __A16_NET_214;
    wire __A16_NET_215;
    wire __A16_NET_216;
    wire __A16_NET_217;
    wire __A16_NET_218;
    wire __A16_NET_219;
    wire __A16_NET_220;
    wire __A16_NET_221;
    wire __A16_NET_222;
    wire __A16_NET_223;
    wire __A16_NET_224;
    wire __A16_NET_225;
    wire __A16_NET_226;
    wire __A16_NET_227;
    wire __A16_NET_228;
    wire __A16_NET_229;
    wire __A16_NET_230;
    wire __A16_NET_231;
    wire __A16_NET_232;
    wire __A16_NET_233;
    wire __A16_NET_234;
    wire __A16_NET_235;
    wire __A16_NET_236;
    wire __A16_NET_237;
    wire __A16_NET_238;
    wire __A16_NET_239;
    wire __A16_NET_240;
    wire __A16_NET_241;
    wire __A16_NET_242;
    wire __A16_NET_243;
    wire __A16_NET_244;
    wire __A16_NET_245;
    wire __A16_NET_246;
    wire __A16_NET_247;
    wire __A16_NET_248;
    wire __A16_NET_249;
    wire __A16_NET_250;
    wire __A16_NET_251;
    wire __A16_NET_252;
    wire __A16_NET_253;
    wire __A16_NET_254;
    wire __A16_NET_255;
    wire __A16_NET_256;
    wire __A16_NET_257;
    wire __A16_NET_258;
    wire __A16_NET_259;
    wire __A16_NET_260;
    wire __A16_NET_261;
    wire __A16_NET_262;
    wire __A16_NET_263;
    wire __A16_NET_264;
    wire __A16_NET_265;
    wire __A16_NET_266;
    wire __A16_NET_267;
    wire __A16_NET_268;
    wire __A16_NET_269;
    wire __A16_NET_270;
    wire __A16_NET_271;
    wire __A16_NET_272;
    wire __A16_NET_273;
    wire __A16_NET_274;
    wire __A16_NET_275;
    wire __A16_NET_276;
    wire __A16_NET_277;
    wire __A16_NET_278;
    wire __A16_NET_279;
    wire __A16_NET_280;
    wire __A16_NET_281;
    wire __A17_1__CH3209;
    wire __A17_1__CH3210;
    wire __A17_1__CH3313;
    wire __A17_1__CH3314;
    wire __A17_1__CH3316;
    wand __A17_1__CHOR01_n;
    wire __A17_1__CHOR01_n_U17004_2;
    wand __A17_1__CHOR02_n;
    wire __A17_1__CHOR02_n_U17004_4;
    wand __A17_1__CHOR03_n;
    wire __A17_1__CHOR03_n_U17004_6;
    wand __A17_1__CHOR04_n;
    wire __A17_1__CHOR04_n_U17004_8;
    wand __A17_1__CHOR05_n;
    wire __A17_1__CHOR05_n_U17004_10;
    wand __A17_1__CHOR06_n;
    wire __A17_1__CHOR06_n_U17004_12;
    wand __A17_1__CHOR07_n;
    wire __A17_1__CHOR07_n_U17013_2;
    wand __A17_1__CHOR08_n;
    wire __A17_1__CHOR08_n_U17013_4;
    wand __A17_1__CHOR09_n;
    wire __A17_1__CHOR09_n_U17013_6;
    wand __A17_1__CHOR10_n;
    wire __A17_1__CHOR10_n_U17013_8;
    wand __A17_1__CHOR11_n;
    wire __A17_1__CHOR11_n_U17013_10;
    wand __A17_1__CHOR12_n;
    wire __A17_1__CHOR12_n_U17013_12;
    wand __A17_1__CHOR13_n;
    wire __A17_1__CHOR13_n_U17020_2;
    wand __A17_1__CHOR14_n;
    wire __A17_1__CHOR14_n_U17020_4;
    wand __A17_1__CHOR16_n;
    wire __A17_1__CHOR16_n_U17020_6;
    wire __A17_1__F04B_n;
    wire __A17_1__FO5D;
    wire __A17_1__HNDRPT;
    wire __A17_1__RCH30_n;
    wire __A17_1__RCH31_n;
    wire __A17_1__RCH32_n;
    wire __A17_1__RCH33_n;
    wire __A17_1__TRP31A;
    wire __A17_1__TRP31B;
    wire __A17_1__TRP32;
    wire __A17_2__CCH10;
    wand __A17_2__CHOR01_n;
    wire __A17_2__CHOR01_n_U17028_10;
    wand __A17_2__CHOR02_n;
    wire __A17_2__CHOR02_n_U17042_2;
    wand __A17_2__CHOR03_n;
    wire __A17_2__CHOR03_n_U17042_4;
    wand __A17_2__CHOR04_n;
    wire __A17_2__CHOR04_n_U17042_6;
    wand __A17_2__CHOR05_n;
    wire __A17_2__CHOR05_n_U17042_8;
    wand __A17_2__CHOR06_n;
    wire __A17_2__CHOR06_n_U17042_10;
    wand __A17_2__CHOR07_n;
    wire __A17_2__CHOR07_n_U17028_12;
    wand __A17_2__CHOR08_n;
    wire __A17_2__CHOR08_n_U17042_12;
    wand __A17_2__CHOR09_n;
    wire __A17_2__CHOR09_n_U17053_2;
    wand __A17_2__CHOR10_n;
    wire __A17_2__CHOR10_n_U17053_4;
    wand __A17_2__CHOR11_n;
    wire __A17_2__CHOR11_n_U17053_6;
    wand __A17_2__CHOR12_n;
    wire __A17_2__CHOR12_n_U17053_8;
    wand __A17_2__CHOR13_n;
    wire __A17_2__CHOR13_n_U17053_10;
    wand __A17_2__CHOR14_n;
    wire __A17_2__CHOR14_n_U17053_12;
    wand __A17_2__CHOR16_n;
    wire __A17_2__CHOR16_n_U17062_2;
    wire __A17_2__RCH10_n;
    wire __A17_2__RLYB01;
    wire __A17_2__RLYB02;
    wire __A17_2__RLYB03;
    wire __A17_2__RLYB04;
    wire __A17_2__RLYB05;
    wire __A17_2__RLYB06;
    wire __A17_2__RLYB07;
    wire __A17_2__RLYB08;
    wire __A17_2__RLYB09;
    wire __A17_2__RLYB10;
    wire __A17_2__RLYB11;
    wire __A17_2__RYWD12;
    wire __A17_2__RYWD13;
    wire __A17_2__RYWD14;
    wire __A17_2__RYWD16;
    wire __A17_2__WCH10_n;
    wire __A17_NET_190;
    wire __A17_NET_191;
    wire __A17_NET_192;
    wire __A17_NET_193;
    wire __A17_NET_194;
    wire __A17_NET_195;
    wire __A17_NET_196;
    wire __A17_NET_197;
    wire __A17_NET_198;
    wire __A17_NET_199;
    wire __A17_NET_200;
    wire __A17_NET_201;
    wire __A17_NET_202;
    wire __A17_NET_203;
    wire __A17_NET_204;
    wire __A17_NET_205;
    wand __A17_NET_207;
    wire __A17_NET_207_U17020_10;
    wire __A17_NET_207_U17020_8;
    wire __A17_NET_208;
    wire __A17_NET_209;
    wire __A17_NET_210;
    wire __A17_NET_211;
    wire __A17_NET_212;
    wire __A17_NET_213;
    wire __A17_NET_214;
    wire __A17_NET_215;
    wire __A17_NET_216;
    wire __A17_NET_217;
    wire __A17_NET_218;
    wire __A17_NET_219;
    wire __A17_NET_220;
    wire __A17_NET_221;
    wire __A17_NET_222;
    wire __A17_NET_223;
    wire __A17_NET_224;
    wire __A17_NET_225;
    wire __A17_NET_226;
    wire __A17_NET_227;
    wire __A17_NET_228;
    wire __A17_NET_229;
    wire __A17_NET_230;
    wire __A17_NET_231;
    wire __A17_NET_232;
    wire __A17_NET_233;
    wire __A17_NET_234;
    wire __A17_NET_235;
    wire __A17_NET_236;
    wire __A17_NET_237;
    wire __A17_NET_238;
    wire __A17_NET_239;
    wire __A17_NET_240;
    wire __A17_NET_241;
    wire __A17_NET_242;
    wire __A17_NET_243;
    wire __A17_NET_244;
    wire __A17_NET_245;
    wire __A17_NET_246;
    wire __A17_NET_247;
    wire __A17_NET_248;
    wire __A17_NET_249;
    wire __A17_NET_250;
    wire __A17_NET_251;
    wire __A17_NET_252;
    wire __A17_NET_253;
    wand __A17_NET_254;
    wire __A17_NET_254_U17020_12;
    wire __A17_NET_254_U17028_2;
    wire __A17_NET_255;
    wire __A17_NET_256;
    wire __A17_NET_257;
    wire __A17_NET_258;
    wire __A17_NET_259;
    wire __A17_NET_261;
    wire __A17_NET_262;
    wire __A17_NET_264;
    wand __A17_NET_265;
    wire __A17_NET_265_U17028_4;
    wire __A17_NET_265_U17028_6;
    wire __A17_NET_265_U17028_8;
    wire __A17_NET_266;
    wire __A17_NET_267;
    wire __A17_NET_268;
    wire __A17_NET_269;
    wire __A17_NET_270;
    wire __A17_NET_271;
    wire __A17_NET_272;
    wire __A17_NET_273;
    wire __A17_NET_274;
    wire __A17_NET_275;
    wire __A17_NET_276;
    wire __A17_NET_277;
    wire __A17_NET_278;
    wire __A17_NET_280;
    wire __A17_NET_281;
    wire __A17_NET_282;
    wire __A17_NET_283;
    wire __A17_NET_284;
    wire __A17_NET_285;
    wire __A17_NET_286;
    wire __A17_NET_287;
    wire __A17_NET_288;
    wire __A17_NET_289;
    wire __A17_NET_290;
    wire __A17_NET_291;
    wire __A17_NET_292;
    wire __A17_NET_293;
    wire __A17_NET_294;
    wire __A17_NET_295;
    wire __A17_NET_296;
    wire __A17_NET_297;
    wire __A17_NET_298;
    wire __A17_NET_299;
    wire __A17_NET_300;
    wire __A17_NET_301;
    wire __A17_NET_302;
    wire __A17_NET_303;
    wire __A17_NET_304;
    wire __A17_NET_305;
    wire __A17_NET_306;
    wire __A17_NET_307;
    wire __A17_NET_308;
    wire __A17_NET_309;
    wire __A17_NET_310;
    wire __A17_NET_311;
    wire __A17_NET_312;
    wire __A17_NET_313;
    wire __A17_NET_314;
    wire __A17_NET_315;
    wire __A17_NET_316;
    wire __A17_NET_317;
    wire __A17_NET_318;
    wire __A17_NET_319;
    wire __A17_NET_320;
    wire __A17_NET_321;
    wire __A17_NET_322;
    wire __A17_NET_323;
    wire __A17_NET_324;
    wire __A17_NET_325;
    wire __A17_NET_326;
    wire __A17_NET_327;
    wire __A17_NET_328;
    wire __A17_NET_329;
    wire __A17_NET_330;
    wire __A17_NET_331;
    wire __A17_NET_332;
    wire __A17_NET_333;
    wire __A17_NET_334;
    wire __A17_NET_336;
    wire __A17_NET_337;
    wire __A17_NET_339;
    wire __A17_NET_340;
    wire __A17_NET_341;
    wire __A17_NET_342;
    wire __A17_NET_343;
    wire __A17_NET_344;
    wire __A17_NET_345;
    wire __A17_NET_346;
    wire __A17_NET_347;
    wire __A17_NET_348;
    wire __A17_NET_349;
    wire __A17_NET_350;
    wire __A17_NET_351;
    wire __A17_NET_352;
    wire __A17_NET_353;
    wire __A17_NET_354;
    wire __A17_NET_355;
    wire __A17_NET_356;
    wire __A17_NET_357;
    wire __A17_NET_358;
    wire __A17_NET_359;
    wire __A17_NET_360;
    wire __A17_NET_361;
    wire __A17_NET_363;
    wire __A17_NET_364;
    wire __A17_NET_365;
    wire __A17_NET_366;
    wire __A17_NET_367;
    wire __A17_NET_368;
    wire __A17_NET_369;
    wire __A17_NET_370;
    wire __A17_NET_371;
    wire __A18_1__CH1505;
    wire __A18_1__CH1601;
    wire __A18_1__CH1602;
    wire __A18_1__CH1603;
    wire __A18_1__CH1604;
    wire __A18_1__CH1605;
    wire __A18_1__CH1606;
    wire __A18_1__CH1607;
    wire __A18_1__F08B_n;
    wire __A18_1__F09A_n;
    wire __A18_1__F09D;
    wire __A18_1__F17A_n;
    wire __A18_1__F17B_n;
    wire __A18_1__RCH15_n;
    wire __A18_1__RCH16_n;
    wire __A18_1__SBYLIT;
    wire __A18_1__STNDBY;
    wire __A18_2__ACTV_n;
    wire __A18_2__ADVCNT;
    wand __A18_2__CNTOF9;
    wire __A18_2__CNTOF9_U18007_10;
    wire __A18_2__CNTOF9_U18007_12;
    wire __A18_2__F10AS0;
    wire __A18_2__HERB;
    wire __A18_2__LRRANG;
    wire __A18_2__LRXVEL;
    wire __A18_2__LRYVEL;
    wire __A18_2__LRZVEL;
    wire __A18_2__RRRANG;
    wire __A18_2__RRRARA;
    wire __A18_NET_100;
    wire __A18_NET_101;
    wire __A18_NET_102;
    wire __A18_NET_103;
    wire __A18_NET_104;
    wire __A18_NET_105;
    wire __A18_NET_106;
    wire __A18_NET_107;
    wire __A18_NET_108;
    wire __A18_NET_109;
    wire __A18_NET_110;
    wand __A18_NET_111;
    wire __A18_NET_111_U18007_2;
    wire __A18_NET_111_U18007_4;
    wire __A18_NET_112;
    wire __A18_NET_113;
    wire __A18_NET_114;
    wire __A18_NET_115;
    wire __A18_NET_116;
    wire __A18_NET_117;
    wire __A18_NET_118;
    wire __A18_NET_119;
    wire __A18_NET_120;
    wire __A18_NET_121;
    wire __A18_NET_122;
    wire __A18_NET_123;
    wire __A18_NET_124;
    wire __A18_NET_125;
    wire __A18_NET_126;
    wire __A18_NET_127;
    wire __A18_NET_128;
    wire __A18_NET_129;
    wire __A18_NET_131;
    wire __A18_NET_134;
    wire __A18_NET_136;
    wire __A18_NET_137;
    wire __A18_NET_138;
    wire __A18_NET_139;
    wire __A18_NET_140;
    wire __A18_NET_141;
    wire __A18_NET_142;
    wire __A18_NET_143;
    wire __A18_NET_144;
    wire __A18_NET_146;
    wire __A18_NET_147;
    wire __A18_NET_148;
    wire __A18_NET_149;
    wire __A18_NET_150;
    wire __A18_NET_151;
    wire __A18_NET_152;
    wand __A18_NET_153;
    wire __A18_NET_153_U18007_6;
    wire __A18_NET_153_U18007_8;
    wire __A18_NET_154;
    wire __A18_NET_155;
    wire __A18_NET_156;
    wire __A18_NET_157;
    wire __A18_NET_158;
    wire __A18_NET_159;
    wire __A18_NET_160;
    wire __A18_NET_161;
    wire __A18_NET_162;
    wire __A18_NET_164;
    wire __A18_NET_165;
    wire __A18_NET_166;
    wire __A18_NET_167;
    wire __A18_NET_168;
    wire __A18_NET_169;
    wire __A18_NET_170;
    wire __A18_NET_172;
    wire __A18_NET_173;
    wire __A18_NET_174;
    wire __A18_NET_175;
    wire __A18_NET_176;
    wire __A18_NET_177;
    wire __A18_NET_178;
    wire __A18_NET_179;
    wire __A18_NET_180;
    wire __A18_NET_184;
    wire __A18_NET_185;
    wire __A18_NET_186;
    wire __A18_NET_190;
    wire __A18_NET_191;
    wire __A18_NET_192;
    wire __A18_NET_193;
    wire __A18_NET_194;
    wire __A18_NET_195;
    wire __A18_NET_196;
    wire __A18_NET_197;
    wire __A18_NET_198;
    wire __A18_NET_199;
    wire __A18_NET_200;
    wire __A18_NET_201;
    wire __A18_NET_202;
    wire __A18_NET_203;
    wire __A18_NET_204;
    wire __A18_NET_205;
    wire __A18_NET_206;
    wire __A18_NET_207;
    wire __A18_NET_208;
    wire __A18_NET_209;
    wire __A18_NET_210;
    wire __A18_NET_211;
    wire __A18_NET_212;
    wire __A18_NET_213;
    wire __A18_NET_214;
    wire __A18_NET_215;
    wire __A18_NET_216;
    wire __A18_NET_217;
    wire __A18_NET_218;
    wire __A18_NET_219;
    wire __A18_NET_220;
    wire __A18_NET_221;
    wire __A18_NET_223;
    wire __A18_NET_224;
    wire __A18_NET_225;
    wire __A18_NET_226;
    wire __A18_NET_228;
    wire __A18_NET_229;
    wire __A18_NET_230;
    wire __A18_NET_231;
    wire __A18_NET_232;
    wire __A18_NET_236;
    wire __A18_NET_237;
    wire __A18_NET_238;
    wire __A18_NET_240;
    wire __A18_NET_241;
    wire __A18_NET_242;
    wire __A18_NET_243;
    wire __A18_NET_244;
    wire __A18_NET_245;
    wire __A18_NET_246;
    wire __A18_NET_247;
    wire __A18_NET_248;
    wire __A18_NET_249;
    wire __A18_NET_250;
    wire __A18_NET_251;
    wire __A18_NET_252;
    wire __A18_NET_257;
    wire __A18_NET_258;
    wire __A18_NET_259;
    wire __A18_NET_260;
    wire __A18_NET_261;
    wire __A18_NET_262;
    wire __A18_NET_263;
    wire __A18_NET_266;
    wire __A18_NET_267;
    wire __A18_NET_268;
    wire __A18_NET_269;
    wire __A18_NET_270;
    wire __A18_NET_89;
    wire __A18_NET_90;
    wire __A18_NET_91;
    wire __A18_NET_92;
    wire __A18_NET_93;
    wire __A18_NET_94;
    wire __A18_NET_95;
    wire __A18_NET_96;
    wire __A18_NET_97;
    wire __A18_NET_98;
    wire __A18_NET_99;
    wire __A19_1__ALRT0;
    wire __A19_1__ALRT1;
    wire __A19_1__ALT0;
    wire __A19_1__ALT1;
    wire __A19_1__ALTSNC;
    wire __A19_1__BLKUPL;
    wire __A19_1__C45R_n;
    wire __A19_1__CH3311;
    wire __A19_1__EMSm;
    wire __A19_1__EMSp;
    wire __A19_1__F5ASB0;
    wire __A19_1__F5ASB0_n;
    wire __A19_1__F5ASB2;
    wire __A19_1__F5BSB2;
    wire __A19_1__OTLNK0;
    wire __A19_1__OTLNK1;
    wire __A19_1__SH3MS_n;
    wire __A19_1__THRSTm;
    wire __A19_1__THRSTp;
    wire __A19_1__UPL0_n;
    wire __A19_1__UPL1_n;
    wire __A19_1__UPRUPT;
    wire __A19_1__XLNK0_n;
    wire __A19_1__XLNK1_n;
    wire __A19_2__CH1109;
    wire __A19_2__CH1110;
    wire __A19_2__CH1111;
    wire __A19_2__CH1112;
    wire __A19_2__CNTRSB_n;
    wire __A19_2__ERRST;
    wire __A19_2__F06B_n;
    wire __A19_2__F07C_n;
    wire __A19_2__F07D_n;
    wire __A19_2__F10B_n;
    wire __A19_2__F7CSB1_n;
    wire __A19_2__FF1109_n;
    wire __A19_2__FF1110_n;
    wire __A19_2__FF1111_n;
    wire __A19_2__FF1112_n;
    wire __A19_2__GYENAB;
    wire __A19_2__GYRRST;
    wire __A19_2__GYRSET;
    wire __A19_2__GYXM;
    wire __A19_2__GYXP;
    wire __A19_2__GYYM;
    wire __A19_2__GYYP;
    wire __A19_2__GYZM;
    wire __A19_2__GYZP;
    wire __A19_2__O44;
    wire __A19_2__OT1110;
    wire __A19_2__OT1111;
    wire __A19_2__OT1112;
    wire __A19_2__OUTCOM;
    wire __A19_2__RHCGO;
    wire __A19_NET_158;
    wire __A19_NET_159;
    wire __A19_NET_160;
    wire __A19_NET_162;
    wire __A19_NET_163;
    wire __A19_NET_164;
    wire __A19_NET_165;
    wire __A19_NET_166;
    wire __A19_NET_167;
    wire __A19_NET_168;
    wire __A19_NET_169;
    wire __A19_NET_170;
    wire __A19_NET_171;
    wire __A19_NET_172;
    wire __A19_NET_173;
    wire __A19_NET_175;
    wire __A19_NET_176;
    wire __A19_NET_178;
    wire __A19_NET_179;
    wire __A19_NET_180;
    wire __A19_NET_181;
    wire __A19_NET_182;
    wire __A19_NET_184;
    wire __A19_NET_185;
    wire __A19_NET_186;
    wire __A19_NET_187;
    wire __A19_NET_188;
    wire __A19_NET_189;
    wire __A19_NET_190;
    wire __A19_NET_191;
    wire __A19_NET_194;
    wire __A19_NET_196;
    wire __A19_NET_197;
    wire __A19_NET_198;
    wire __A19_NET_199;
    wire __A19_NET_200;
    wire __A19_NET_201;
    wire __A19_NET_202;
    wire __A19_NET_203;
    wire __A19_NET_204;
    wire __A19_NET_205;
    wire __A19_NET_206;
    wire __A19_NET_207;
    wire __A19_NET_208;
    wire __A19_NET_209;
    wire __A19_NET_210;
    wire __A19_NET_211;
    wire __A19_NET_212;
    wire __A19_NET_213;
    wire __A19_NET_214;
    wire __A19_NET_215;
    wire __A19_NET_216;
    wire __A19_NET_217;
    wire __A19_NET_218;
    wire __A19_NET_219;
    wire __A19_NET_220;
    wire __A19_NET_221;
    wire __A19_NET_222;
    wire __A19_NET_223;
    wire __A19_NET_224;
    wire __A19_NET_225;
    wire __A19_NET_226;
    wire __A19_NET_227;
    wire __A19_NET_228;
    wire __A19_NET_229;
    wire __A19_NET_230;
    wire __A19_NET_231;
    wire __A19_NET_232;
    wire __A19_NET_234;
    wire __A19_NET_235;
    wire __A19_NET_236;
    wire __A19_NET_238;
    wire __A19_NET_239;
    wire __A19_NET_240;
    wire __A19_NET_241;
    wire __A19_NET_242;
    wire __A19_NET_243;
    wire __A19_NET_244;
    wire __A19_NET_245;
    wire __A19_NET_246;
    wire __A19_NET_247;
    wire __A19_NET_248;
    wire __A19_NET_249;
    wire __A19_NET_250;
    wire __A19_NET_251;
    wire __A19_NET_252;
    wire __A19_NET_253;
    wire __A19_NET_254;
    wire __A19_NET_255;
    wire __A19_NET_256;
    wire __A19_NET_257;
    wire __A19_NET_258;
    wire __A19_NET_259;
    wire __A19_NET_260;
    wire __A19_NET_261;
    wire __A19_NET_262;
    wire __A19_NET_263;
    wire __A19_NET_264;
    wire __A19_NET_265;
    wire __A19_NET_266;
    wire __A19_NET_267;
    wire __A19_NET_268;
    wire __A19_NET_269;
    wire __A19_NET_270;
    wire __A19_NET_271;
    wire __A19_NET_272;
    wire __A19_NET_273;
    wire __A19_NET_274;
    wire __A19_NET_275;
    wire __A19_NET_276;
    wire __A19_NET_277;
    wire __A19_NET_278;
    wire __A19_NET_279;
    wire __A19_NET_280;
    wire __A19_NET_281;
    wire __A19_NET_282;
    wire __A19_NET_283;
    wire __A19_NET_284;
    wire __A19_NET_285;
    wire __A19_NET_286;
    wire __A19_NET_287;
    wire __A19_NET_288;
    wire __A19_NET_289;
    wire __A19_NET_290;
    wire __A19_NET_291;
    wire __A19_NET_292;
    wire __A19_NET_293;
    wire __A19_NET_294;
    wire __A19_NET_295;
    wire __A19_NET_296;
    wire __A19_NET_297;
    wire __A19_NET_298;
    wire __A19_NET_299;
    wire __A19_NET_300;
    wire __A19_NET_302;
    wire __A19_NET_303;
    wire __A19_NET_304;
    wire __A19_NET_305;
    wire __A19_NET_311;
    wire __A19_NET_312;
    wire __A19_NET_313;
    wire __A19_NET_314;
    wire __A19_NET_315;
    wire __A19_NET_316;
    wire __A19_NET_317;
    wire __A19_NET_318;
    wire __A19_NET_319;
    wire __A19_NET_320;
    wire __A19_NET_321;
    wire __A19_NET_322;
    wire __A19_NET_323;
    wire __A19_NET_324;
    wire __A19_NET_325;
    wire __A19_NET_326;
    wire __A20_1__C10R;
    wire __A20_1__C1R;
    wire __A20_1__C2R;
    wire __A20_1__C3R;
    wire __A20_1__C4R;
    wire __A20_1__C5R;
    wire __A20_1__C6R;
    wire __A20_1__C7R;
    wire __A20_1__C8R;
    wire __A20_1__C9R;
    wire __A20_1___CG1;
    wire __A20_1___CG2OUT;
    wire __A20_1___CG5OUT;
    wire __A20_2__C10R;
    wire __A20_2__C1R;
    wire __A20_2__C2R;
    wire __A20_2__C3R;
    wire __A20_2__C4R;
    wire __A20_2__C5R;
    wire __A20_2__C6R;
    wire __A20_2__C7R;
    wire __A20_2__C8R;
    wire __A20_2__C9R;
    wire __A20_2___CG1;
    wire __A20_2___CG10OUT;
    wire __A20_2___CG6;
    wire __A20_NET_100;
    wire __A20_NET_101;
    wire __A20_NET_102;
    wire __A20_NET_103;
    wire __A20_NET_104;
    wire __A20_NET_106;
    wire __A20_NET_107;
    wire __A20_NET_108;
    wire __A20_NET_109;
    wire __A20_NET_111;
    wire __A20_NET_112;
    wire __A20_NET_115;
    wire __A20_NET_118;
    wire __A20_NET_119;
    wire __A20_NET_120;
    wire __A20_NET_121;
    wire __A20_NET_122;
    wire __A20_NET_124;
    wire __A20_NET_125;
    wire __A20_NET_126;
    wire __A20_NET_127;
    wire __A20_NET_128;
    wire __A20_NET_129;
    wire __A20_NET_131;
    wire __A20_NET_132;
    wire __A20_NET_133;
    wire __A20_NET_134;
    wire __A20_NET_135;
    wire __A20_NET_136;
    wire __A20_NET_137;
    wire __A20_NET_138;
    wire __A20_NET_139;
    wire __A20_NET_140;
    wire __A20_NET_141;
    wire __A20_NET_142;
    wire __A20_NET_144;
    wire __A20_NET_145;
    wire __A20_NET_146;
    wire __A20_NET_147;
    wire __A20_NET_148;
    wire __A20_NET_150;
    wire __A20_NET_151;
    wire __A20_NET_152;
    wire __A20_NET_153;
    wire __A20_NET_154;
    wire __A20_NET_156;
    wire __A20_NET_157;
    wire __A20_NET_162;
    wire __A20_NET_163;
    wire __A20_NET_164;
    wire __A20_NET_165;
    wire __A20_NET_166;
    wire __A20_NET_167;
    wire __A20_NET_168;
    wire __A20_NET_169;
    wire __A20_NET_170;
    wire __A20_NET_172;
    wire __A20_NET_173;
    wire __A20_NET_174;
    wire __A20_NET_176;
    wire __A20_NET_177;
    wire __A20_NET_178;
    wire __A20_NET_179;
    wire __A20_NET_180;
    wire __A20_NET_181;
    wire __A20_NET_182;
    wire __A20_NET_183;
    wire __A20_NET_184;
    wire __A20_NET_185;
    wire __A20_NET_186;
    wire __A20_NET_188;
    wire __A20_NET_189;
    wire __A20_NET_190;
    wire __A20_NET_191;
    wire __A20_NET_192;
    wire __A20_NET_194;
    wire __A20_NET_195;
    wire __A20_NET_196;
    wire __A20_NET_197;
    wire __A20_NET_199;
    wire __A20_NET_200;
    wire __A20_NET_203;
    wire __A20_NET_206;
    wire __A20_NET_207;
    wire __A20_NET_208;
    wire __A20_NET_209;
    wire __A20_NET_210;
    wire __A20_NET_212;
    wire __A20_NET_213;
    wire __A20_NET_214;
    wire __A20_NET_215;
    wire __A20_NET_216;
    wire __A20_NET_217;
    wire __A20_NET_219;
    wire __A20_NET_220;
    wire __A20_NET_221;
    wire __A20_NET_222;
    wire __A20_NET_223;
    wire __A20_NET_224;
    wire __A20_NET_225;
    wire __A20_NET_226;
    wire __A20_NET_227;
    wire __A20_NET_228;
    wire __A20_NET_229;
    wire __A20_NET_230;
    wire __A20_NET_232;
    wire __A20_NET_233;
    wire __A20_NET_234;
    wire __A20_NET_235;
    wire __A20_NET_236;
    wire __A20_NET_238;
    wire __A20_NET_239;
    wire __A20_NET_240;
    wire __A20_NET_241;
    wire __A20_NET_243;
    wire __A20_NET_244;
    wire __A20_NET_246;
    wire __A20_NET_250;
    wire __A20_NET_251;
    wire __A20_NET_252;
    wire __A20_NET_253;
    wire __A20_NET_254;
    wire __A20_NET_256;
    wire __A20_NET_257;
    wire __A20_NET_258;
    wire __A20_NET_259;
    wire __A20_NET_261;
    wire __A20_NET_262;
    wire __A20_NET_263;
    wire __A20_NET_264;
    wire __A20_NET_265;
    wire __A20_NET_90;
    wire __A20_NET_91;
    wire __A20_NET_92;
    wire __A20_NET_93;
    wire __A20_NET_94;
    wire __A20_NET_95;
    wire __A20_NET_96;
    wire __A20_NET_97;
    wire __A20_NET_98;
    wire __A21_1__30SUM;
    wand __A21_1__32004K;
    wire __A21_1__32004K_U21010_2;
    wire __A21_1__32004K_U21010_4;
    wire __A21_1__50SUM;
    wire __A21_1__C42A;
    wire __A21_1__C42M;
    wire __A21_1__C42P;
    wire __A21_1__C43A;
    wire __A21_1__C43M;
    wire __A21_1__C43P;
    wire __A21_1__C44A;
    wire __A21_1__C44M;
    wire __A21_1__C44P;
    wire __A21_1__C45A;
    wire __A21_1__C45M;
    wire __A21_1__C45P;
    wire __A21_1__C46A;
    wire __A21_1__C46M;
    wire __A21_1__C46P;
    wire __A21_1__C47A;
    wire __A21_1__C56A;
    wire __A21_1__C57A;
    wire __A21_1__C60A;
    wire __A21_1__DINCNC_n;
    wire __A21_1__MCDU_n;
    wire __A21_1__MINC_n;
    wire __A21_1__PCDU_n;
    wire __A21_1__PINC_n;
    wire __A21_1__RSCT_n;
    wire __A21_1__SHANC;
    wire __A21_1__SHINC;
    wire __A21_3__C42R;
    wire __A21_3__C43R;
    wire __A21_3__C44R;
    wire __A21_3__C46R;
    wire __A21_3__C47R;
    wire __A21_3__C56R;
    wire __A21_3__C57R;
    wire __A21_3__C60R;
    wire __A21_3__CG15;
    wire __A21_3__CG16;
    wire __A21_NET_132;
    wand __A21_NET_133;
    wire __A21_NET_133_U21024_2;
    wire __A21_NET_133_U21024_4;
    wire __A21_NET_133_U21024_6;
    wire __A21_NET_134;
    wire __A21_NET_138;
    wire __A21_NET_140;
    wire __A21_NET_141;
    wand __A21_NET_142;
    wire __A21_NET_142_U21024_10;
    wire __A21_NET_142_U21024_8;
    wire __A21_NET_143;
    wire __A21_NET_144;
    wand __A21_NET_145;
    wire __A21_NET_145_U21010_10;
    wire __A21_NET_145_U21010_12;
    wand __A21_NET_146;
    wire __A21_NET_146_U21006_10;
    wire __A21_NET_146_U21006_12;
    wire __A21_NET_146_U21006_6;
    wire __A21_NET_146_U21006_8;
    wand __A21_NET_147;
    wire __A21_NET_147_U21002_10;
    wire __A21_NET_147_U21002_12;
    wire __A21_NET_147_U21006_2;
    wire __A21_NET_147_U21006_4;
    wire __A21_NET_148;
    wand __A21_NET_149;
    wire __A21_NET_149_U21010_6;
    wire __A21_NET_149_U21010_8;
    wire __A21_NET_150;
    wire __A21_NET_152;
    wire __A21_NET_153;
    wire __A21_NET_154;
    wire __A21_NET_155;
    wand __A21_NET_157;
    wire __A21_NET_157_U21024_12;
    wire __A21_NET_157_U21028_2;
    wire __A21_NET_158;
    wand __A21_NET_159;
    wire __A21_NET_159_U21028_4;
    wire __A21_NET_159_U21028_6;
    wire __A21_NET_160;
    wire __A21_NET_161;
    wire __A21_NET_162;
    wire __A21_NET_163;
    wire __A21_NET_164;
    wire __A21_NET_167;
    wire __A21_NET_168;
    wire __A21_NET_169;
    wire __A21_NET_172;
    wire __A21_NET_173;
    wire __A21_NET_182;
    wire __A21_NET_183;
    wire __A21_NET_184;
    wire __A21_NET_189;
    wire __A21_NET_193;
    wire __A21_NET_198;
    wire __A21_NET_203;
    wire __A21_NET_204;
    wand __A21_NET_205;
    wire __A21_NET_205_U21002_2;
    wire __A21_NET_205_U21002_4;
    wire __A21_NET_205_U21002_6;
    wire __A21_NET_205_U21002_8;
    wire __A21_NET_206;
    wire __A21_NET_207;
    wire __A21_NET_209;
    wire __A21_NET_211;
    wire __A21_NET_212;
    wire __A21_NET_217;
    wire __A21_NET_220;
    wire __A21_NET_221;
    wire __A21_NET_222;
    wand __A21_NET_223;
    wire __A21_NET_223_U21015_2;
    wire __A21_NET_223_U21015_4;
    wire __A21_NET_223_U21015_6;
    wire __A21_NET_228;
    wand __A21_NET_229;
    wire __A21_NET_229_U21015_10;
    wire __A21_NET_229_U21015_12;
    wire __A21_NET_229_U21015_8;
    wire __A21_NET_230;
    wire __A21_NET_231;
    wire __A21_NET_232;
    wire __A21_NET_233;
    wire __A21_NET_234;
    wire __A21_NET_235;
    wire __A21_NET_237;
    wire __A21_NET_238;
    wire __A21_NET_239;
    wire __A21_NET_240;
    wire __A21_NET_241;
    wire __A21_NET_242;
    wire __A21_NET_243;
    wire __A21_NET_244;
    wire __A21_NET_245;
    wire __A21_NET_246;
    wire __A21_NET_247;
    wire __A21_NET_248;
    wire __A21_NET_249;
    wire __A21_NET_250;
    wire __A21_NET_251;
    wire __A21_NET_252;
    wire __A21_NET_253;
    wire __A21_NET_254;
    wire __A21_NET_255;
    wire __A21_NET_256;
    wire __A21_NET_257;
    wire __A21_NET_258;
    wire __A21_NET_259;
    wire __A21_NET_261;
    wire __A21_NET_262;
    wire __A21_NET_263;
    wire __A21_NET_264;
    wire __A21_NET_265;
    wire __A21_NET_266;
    wire __A21_NET_267;
    wire __A21_NET_268;
    wire __A21_NET_269;
    wire __A21_NET_270;
    wire __A21_NET_271;
    wire __A21_NET_272;
    wire __A21_NET_273;
    wire __A21_NET_275;
    wire __A21_NET_276;
    wire __A21_NET_277;
    wire __A21_NET_278;
    wire __A21_NET_279;
    wire __A21_NET_280;
    wire __A21_NET_281;
    wire __A21_NET_282;
    wire __A21_NET_283;
    wire __A21_NET_284;
    wire __A21_NET_285;
    wire __A21_NET_286;
    wire __A21_NET_287;
    wire __A21_NET_288;
    wire __A21_NET_289;
    wire __A21_NET_290;
    wire __A21_NET_291;
    wire __A21_NET_292;
    wire __A21_NET_293;
    wire __A21_NET_294;
    wire __A21_NET_295;
    wire __A21_NET_296;
    wire __A21_NET_297;
    wire __A21_NET_298;
    wire __A21_NET_299;
    wire __A21_NET_300;
    wire __A22_1__16CNT;
    wire __A22_1__1CNT;
    wire __A22_1__32CNT;
    wire __A22_1__ADVCTR;
    wire __A22_1__BSYNC_n;
    wand __A22_1__DATA_n;
    wire __A22_1__DATA_n_U22028_10;
    wire __A22_1__DATA_n_U22028_12;
    wire __A22_1__DATA_n_U22028_2;
    wire __A22_1__DATA_n_U22028_4;
    wire __A22_1__DATA_n_U22028_6;
    wire __A22_1__DATA_n_U22028_8;
    wire __A22_1__DATA_n_U22057_2;
    wire __A22_1__DATA_n_U22057_4;
    wire __A22_1__DKCTR1;
    wire __A22_1__DKCTR1_n;
    wire __A22_1__DKCTR2;
    wire __A22_1__DKCTR2_n;
    wire __A22_1__DKCTR3;
    wire __A22_1__DKCTR3_n;
    wire __A22_1__DKCTR4;
    wire __A22_1__DKCTR4_n;
    wire __A22_1__DKCTR5;
    wire __A22_1__DKCTR5_n;
    wire __A22_1__DKDATA;
    wire __A22_1__DKDATB;
    wire __A22_1__DKDAT_n;
    wire __A22_1__DLKCLR;
    wire __A22_1__DLKRPT;
    wire __A22_1__END;
    wire __A22_1__HIGH0_n;
    wire __A22_1__HIGH1_n;
    wire __A22_1__HIGH2_n;
    wire __A22_1__HIGH3_n;
    wire __A22_1__LOW0_n;
    wire __A22_1__LOW1_n;
    wire __A22_1__LOW2_n;
    wire __A22_1__LOW3_n;
    wire __A22_1__LOW4_n;
    wire __A22_1__LOW5_n;
    wire __A22_1__LOW6_n;
    wire __A22_1__LOW7_n;
    wire __A22_1__ORDRBT;
    wire __A22_1__RDOUT_n;
    wire __A22_1__WDORDR;
    wire __A22_1__WRD1B1;
    wire __A22_1__WRD1BP;
    wire __A22_1__WRD2B2;
    wire __A22_1__WRD2B3;
    wire __A22_NET_101;
    wire __A22_NET_102;
    wire __A22_NET_103;
    wire __A22_NET_104;
    wire __A22_NET_107;
    wire __A22_NET_108;
    wire __A22_NET_109;
    wire __A22_NET_111;
    wire __A22_NET_113;
    wire __A22_NET_114;
    wire __A22_NET_116;
    wire __A22_NET_117;
    wire __A22_NET_118;
    wire __A22_NET_119;
    wire __A22_NET_120;
    wire __A22_NET_121;
    wire __A22_NET_122;
    wire __A22_NET_123;
    wire __A22_NET_124;
    wire __A22_NET_125;
    wire __A22_NET_126;
    wire __A22_NET_127;
    wire __A22_NET_128;
    wire __A22_NET_129;
    wire __A22_NET_130;
    wire __A22_NET_132;
    wire __A22_NET_133;
    wire __A22_NET_134;
    wire __A22_NET_135;
    wire __A22_NET_137;
    wire __A22_NET_138;
    wire __A22_NET_139;
    wire __A22_NET_140;
    wire __A22_NET_141;
    wire __A22_NET_142;
    wire __A22_NET_143;
    wire __A22_NET_144;
    wire __A22_NET_145;
    wire __A22_NET_146;
    wire __A22_NET_147;
    wire __A22_NET_148;
    wire __A22_NET_149;
    wire __A22_NET_150;
    wire __A22_NET_151;
    wire __A22_NET_152;
    wire __A22_NET_153;
    wire __A22_NET_154;
    wire __A22_NET_155;
    wire __A22_NET_156;
    wire __A22_NET_157;
    wire __A22_NET_158;
    wire __A22_NET_159;
    wire __A22_NET_160;
    wire __A22_NET_161;
    wire __A22_NET_162;
    wire __A22_NET_163;
    wire __A22_NET_164;
    wire __A22_NET_165;
    wire __A22_NET_166;
    wire __A22_NET_167;
    wire __A22_NET_168;
    wire __A22_NET_169;
    wire __A22_NET_170;
    wire __A22_NET_171;
    wire __A22_NET_172;
    wire __A22_NET_173;
    wire __A22_NET_174;
    wire __A22_NET_176;
    wire __A22_NET_178;
    wire __A22_NET_179;
    wire __A22_NET_180;
    wire __A22_NET_181;
    wire __A22_NET_182;
    wire __A22_NET_183;
    wire __A22_NET_184;
    wire __A22_NET_185;
    wire __A22_NET_186;
    wire __A22_NET_187;
    wire __A22_NET_190;
    wire __A22_NET_191;
    wire __A22_NET_192;
    wire __A22_NET_193;
    wire __A22_NET_194;
    wire __A22_NET_195;
    wire __A22_NET_196;
    wire __A22_NET_197;
    wire __A22_NET_198;
    wire __A22_NET_199;
    wire __A22_NET_200;
    wire __A22_NET_201;
    wire __A22_NET_202;
    wire __A22_NET_203;
    wire __A22_NET_204;
    wire __A22_NET_207;
    wire __A22_NET_208;
    wire __A22_NET_209;
    wire __A22_NET_210;
    wire __A22_NET_211;
    wire __A22_NET_212;
    wire __A22_NET_213;
    wire __A22_NET_214;
    wire __A22_NET_215;
    wire __A22_NET_216;
    wire __A22_NET_217;
    wire __A22_NET_218;
    wire __A22_NET_219;
    wire __A22_NET_220;
    wire __A22_NET_221;
    wire __A22_NET_222;
    wire __A22_NET_223;
    wire __A22_NET_224;
    wire __A22_NET_225;
    wire __A22_NET_226;
    wire __A22_NET_227;
    wire __A22_NET_228;
    wire __A22_NET_229;
    wire __A22_NET_230;
    wire __A22_NET_231;
    wire __A22_NET_232;
    wire __A22_NET_233;
    wire __A22_NET_234;
    wire __A22_NET_235;
    wire __A22_NET_236;
    wire __A22_NET_239;
    wire __A22_NET_240;
    wire __A22_NET_241;
    wire __A22_NET_242;
    wire __A22_NET_243;
    wire __A22_NET_244;
    wire __A22_NET_246;
    wire __A22_NET_247;
    wire __A22_NET_248;
    wire __A22_NET_249;
    wire __A22_NET_251;
    wire __A22_NET_252;
    wire __A22_NET_253;
    wire __A22_NET_254;
    wire __A22_NET_255;
    wire __A22_NET_256;
    wire __A22_NET_257;
    wire __A22_NET_258;
    wire __A22_NET_259;
    wire __A22_NET_260;
    wire __A22_NET_261;
    wire __A22_NET_262;
    wire __A22_NET_263;
    wire __A22_NET_264;
    wire __A22_NET_265;
    wire __A22_NET_266;
    wire __A22_NET_267;
    wire __A22_NET_268;
    wire __A22_NET_271;
    wire __A22_NET_272;
    wire __A22_NET_273;
    wire __A22_NET_274;
    wire __A22_NET_275;
    wire __A22_NET_276;
    wire __A22_NET_277;
    wire __A22_NET_57;
    wire __A22_NET_58;
    wire __A22_NET_61;
    wire __A22_NET_62;
    wire __A22_NET_63;
    wire __A22_NET_65;
    wire __A22_NET_66;
    wire __A22_NET_67;
    wire __A22_NET_69;
    wire __A22_NET_71;
    wire __A22_NET_72;
    wire __A22_NET_75;
    wire __A22_NET_77;
    wire __A22_NET_78;
    wire __A22_NET_79;
    wire __A22_NET_80;
    wire __A22_NET_81;
    wire __A22_NET_82;
    wire __A22_NET_83;
    wire __A22_NET_84;
    wire __A22_NET_85;
    wire __A22_NET_86;
    wire __A22_NET_87;
    wire __A22_NET_88;
    wire __A22_NET_89;
    wire __A22_NET_90;
    wire __A22_NET_93;
    wire __A22_NET_97;
    wire __A22_NET_98;
    wire __B01_1__CQA;
    wire __B01_1__CQB;
    wire __B01_1__CQC;
    wire __B01_1__FADDR1;
    wire __B01_1__FADDR10;
    wire __B01_1__FADDR11;
    wire __B01_1__FADDR12;
    wire __B01_1__FADDR13;
    wire __B01_1__FADDR14;
    wire __B01_1__FADDR15;
    wire __B01_1__FADDR16;
    wire __B01_1__FADDR2;
    wire __B01_1__FADDR3;
    wire __B01_1__FADDR4;
    wire __B01_1__FADDR5;
    wire __B01_1__FADDR6;
    wire __B01_1__FADDR7;
    wire __B01_1__FADDR8;
    wire __B01_1__FADDR9;
    wire __B01_1__QUARTERA;
    wire __B01_1__QUARTERB;
    wire __B01_1__QUARTERC;
    wire __B01_2__ES01_n;
    wire __B01_2__ES02_n;
    wire __B01_2__ES03_n;
    wire __B01_2__ES04_n;
    wire __B01_2__ES05_n;
    wire __B01_2__ES06_n;
    wire __B01_2__ES07_n;
    wire __B01_2__ES08_n;
    wire __B01_2__ES09_n;
    wire __B01_2__ES10_n;
    wire __B01_2__ES11_n;
    wire __B01_2__RADDR1;
    wire __B01_2__RADDR10;
    wire __B01_2__RADDR11;
    wire __B01_2__RADDR2;
    wire __B01_2__RADDR3;
    wire __B01_2__RADDR4;
    wire __B01_2__RADDR5;
    wire __B01_2__RADDR6;
    wire __B01_2__RADDR7;
    wire __B01_2__RADDR8;
    wire __B01_2__RADDR9;
    wire __B01_2__RESETK;
    wire __B01_NET_101;
    wire __B01_NET_102;
    wire __B01_NET_103;
    wire __B01_NET_104;
    wire __B01_NET_105;
    wire __B01_NET_106;
    wire __B01_NET_108;
    wire __B01_NET_115;
    wire __B01_NET_116;
    wire __B01_NET_118;
    wire __B01_NET_119;
    wire __B01_NET_120;
    wire __B01_NET_121;
    wire __B01_NET_122;
    wire __B01_NET_123;
    wire __B01_NET_124;
    wire __B01_NET_125;
    wire __B01_NET_126;
    wire __B01_NET_128;
    wire __B01_NET_129;
    wire __B01_NET_130;
    wire __B01_NET_131;
    wire __B01_NET_132;
    wire __B01_NET_134;
    wire __B01_NET_135;
    wire __B01_NET_137;
    wire __B01_NET_138;
    wire __B01_NET_139;
    wire __B01_NET_140;
    wire __B01_NET_141;
    wire __B01_NET_142;
    wire __B01_NET_144;
    wire __B01_NET_147;
    wire __B01_NET_148;
    wire __B01_NET_149;
    wire __B01_NET_150;
    wire __B01_NET_155;
    wire __B01_NET_171;
    wire __B01_NET_172;
    wire __B01_NET_173;
    wire __B01_NET_174;
    wire __B01_NET_175;
    wire __B01_NET_176;
    wire __B01_NET_177;
    wire __B01_NET_180;
    wire __B01_NET_181;
    wire __B01_NET_182;
    wire __B01_NET_184;
    wire __B01_NET_185;
    wire __B01_NET_186;
    wire __B01_NET_187;
    wire __B01_NET_188;
    wire __B01_NET_189;
    wire __B01_NET_190;
    wire __B01_NET_192;
    wire __B01_NET_197;
    wire __B01_NET_198;
    wire __B01_NET_200;
    wire __B01_NET_201;
    wire __B01_NET_203;
    wire __B01_NET_204;
    wire __B01_NET_205;
    wire __B01_NET_214;
    wire __B01_NET_215;
    wire __B01_NET_216;
    wire __B01_NET_217;
    wire __B01_NET_218;
    wire __B01_NET_219;
    wire __B01_NET_220;
    wire __B01_NET_221;
    wire __B01_NET_222;
    wire __B01_NET_223;
    wire __B01_NET_224;
    wire __B01_NET_225;
    wire __B01_NET_227;
    wire __B01_NET_230;
    wire __B01_NET_232;
    wire __B01_NET_233;
    wire __B01_NET_235;
    wire __B01_NET_237;
    wire __B01_NET_238;
    wire __B01_NET_239;
    wire __B01_NET_240;
    wire __B01_NET_242;
    wire __B01_NET_243;
    wire __B01_NET_244;
    wire __B01_NET_91;
    wire __B01_NET_92;
    wire __B01_NET_93;
    wire __B01_NET_94;
    wire __B01_NET_96;
    wire __B01_NET_97;
    wire __B01_NET_98;
    wire __B01_NET_99;
    wire n10XP1;
    wire n10XP8;
    wire n11XP2;
    wire n1XP10;
    wire n2XP3;
    wire n2XP5;
    wire n2XP7;
    wire n2XP8;
    wire n3XP2;
    wire n3XP6;
    wire n3XP7;
    wire n4XP11;
    wire n4XP5;
    wand n5XP11;
    wire n5XP11_U4039_6;
    wire n5XP11_U4039_8;
    wire n5XP12;
    wire n5XP15;
    wire n5XP21;
    wire n5XP28;
    wire n5XP4;
    wire n6XP5;
    wire n6XP8;
    wire n7XP14;
    wire n7XP19;
    wire n7XP4;
    wire n7XP9;
    wand n8PP4;
    wire n8PP4_U4063_12;
    wire n8PP4_U6037_10;
    wire n8PP4_U6037_12;
    wire n8PP4_U6041_2;
    wire n8XP5;
    wire n8XP6;
    wire n9XP1;
    wire n9XP5;

    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1001(__A01_1__F02A, __A01_1__scaler_s2__FS_n, __A01_NET_178, __A01_1__F02B, __A01_NET_177, __A01_1__FS02, GND, __A01_NET_178, __A01_1__FS02, __A01_1__scaler_s2__FS_n, __A01_1__scaler_s2__FS_n, __A01_NET_177, __A01_1__FS02, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1002(__A01_1__F02A, FS01_n, __A01_NET_178, FS01_n, __A01_1__F02B, __A01_NET_177, GND, __A01_NET_180, __A01_1__F03A, __A01_1__F02A, __A01_NET_179, __A01_NET_178, __A01_NET_177, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1003(__A01_1__F03A, __A01_1__scaler_s3__FS_n, __A01_NET_180, __A01_1__F03B, __A01_NET_179, __A01_1__FS03, GND, __A01_NET_180, __A01_1__FS03, __A01_1__scaler_s3__FS_n, __A01_1__scaler_s3__FS_n, __A01_NET_179, __A01_1__FS03, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1004(__A01_NET_180, __A01_1__F02A, F04A, __A01_1__F03A, __A01_NET_182, __A01_NET_181, GND, __A01_NET_182, __A01_NET_181, __A01_1__F03A, F04B, __A01_NET_179, __A01_1__F03B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1005(F04A, __A01_1__scaler_s4__FS_n, __A01_NET_181, F04B, __A01_NET_182, __A01_1__FS04, GND, __A01_NET_181, __A01_1__FS04, __A01_1__scaler_s4__FS_n, __A01_1__scaler_s4__FS_n, __A01_NET_182, __A01_1__FS04, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1006(__A01_1__F05A, __A01_1__scaler_s5__FS_n, __A01_NET_184, __A01_1__F05B, __A01_NET_183, __A01_1__FS05, GND, __A01_NET_184, __A01_1__FS05, __A01_1__scaler_s5__FS_n, __A01_1__scaler_s5__FS_n, __A01_NET_183, __A01_1__FS05, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1007(__A01_1__F05A, F04A, __A01_NET_184, F04A, __A01_1__F05B, __A01_NET_183, GND, __A01_NET_185, __A01_1__F06A, __A01_1__F05A, __A01_NET_186, __A01_NET_184, __A01_NET_183, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1008(__A01_1__F06A, __A01_1__scaler_s6__FS_n, __A01_NET_185, F06B, __A01_NET_186, __A01_1__FS06, GND, __A01_NET_185, __A01_1__FS06, __A01_1__scaler_s6__FS_n, __A01_1__scaler_s6__FS_n, __A01_NET_186, __A01_1__FS06, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1009(__A01_NET_185, __A01_1__F05A, F07A, __A01_1__F06A, __A01_NET_187, __A01_NET_188, GND, __A01_NET_187, __A01_NET_188, __A01_1__F06A, F07B, __A01_NET_186, F06B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1010(F07A, __A01_1__scaler_s7__FS_n, __A01_NET_188, F07B, __A01_NET_187, __A01_1__FS07, GND, __A01_NET_188, __A01_1__FS07, __A01_1__scaler_s7__FS_n, __A01_1__scaler_s7__FS_n, __A01_NET_187, __A01_1__FS07, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1011(__A01_1__F08A, __A01_1__scaler_s8__FS_n, __A01_NET_190, F08B, __A01_NET_189, __A01_1__FS08, GND, __A01_NET_190, __A01_1__FS08, __A01_1__scaler_s8__FS_n, __A01_1__scaler_s8__FS_n, __A01_NET_189, __A01_1__FS08, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1012(__A01_1__F08A, F07A, __A01_NET_190, F07A, F08B, __A01_NET_189, GND, __A01_NET_192, F09A, __A01_1__F08A, __A01_NET_191, __A01_NET_190, __A01_NET_189, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1013(F09A, __A01_1__scaler_s9__FS_n, __A01_NET_192, F09B, __A01_NET_191, FS09, GND, __A01_NET_192, FS09, __A01_1__scaler_s9__FS_n, __A01_1__scaler_s9__FS_n, __A01_NET_191, FS09, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1014(__A01_NET_192, __A01_1__F08A, F10A, F09A, __A01_NET_193, __A01_NET_194, GND, __A01_NET_193, __A01_NET_194, F09A, F10B, __A01_NET_191, F09B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1015(F10A, __A01_1__scaler_s10__FS_n, __A01_NET_194, F10B, __A01_NET_193, FS10, GND, __A01_NET_194, FS10, __A01_1__scaler_s10__FS_n, __A01_1__scaler_s10__FS_n, __A01_NET_193, FS10, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1016(__A01_1__F11A, __A01_1__scaler_s11__FS_n, __A01_NET_196, __A01_1__F11B, __A01_NET_195, __A01_1__FS11, GND, __A01_NET_196, __A01_1__FS11, __A01_1__scaler_s11__FS_n, __A01_1__scaler_s11__FS_n, __A01_NET_195, __A01_1__FS11, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1017(__A01_1__F11A, F10A, __A01_NET_196, F10A, __A01_1__F11B, __A01_NET_195, GND, __A01_NET_198, __A01_1__F12A, __A01_1__F11A, __A01_NET_197, __A01_NET_196, __A01_NET_195, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1018(__A01_1__F12A, __A01_1__scaler_s12__FS_n, __A01_NET_198, F12B, __A01_NET_197, __A01_1__FS12, GND, __A01_NET_198, __A01_1__FS12, __A01_1__scaler_s12__FS_n, __A01_1__scaler_s12__FS_n, __A01_NET_197, __A01_1__FS12, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1019(__A01_NET_198, __A01_1__F11A, __A01_1__F13A, __A01_1__F12A, __A01_NET_199, __A01_NET_200, GND, __A01_NET_199, __A01_NET_200, __A01_1__F12A, __A01_1__F13B, __A01_NET_197, F12B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1020(__A01_1__F13A, __A01_1__scaler_s13__FS_n, __A01_NET_200, __A01_1__F13B, __A01_NET_199, FS13, GND, __A01_NET_200, FS13, __A01_1__scaler_s13__FS_n, __A01_1__scaler_s13__FS_n, __A01_NET_199, FS13, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1021(__A01_1__F14A, __A01_1__scaler_s14__FS_n, __A01_NET_201, F14B, __A01_NET_202, FS14, GND, __A01_NET_201, FS14, __A01_1__scaler_s14__FS_n, __A01_1__scaler_s14__FS_n, __A01_NET_202, FS14, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1022(__A01_1__F14A, __A01_1__F13A, __A01_NET_201, __A01_1__F13A, F14B, __A01_NET_202, GND, __A01_NET_204, __A01_1__F15A, __A01_1__F14A, __A01_NET_203, __A01_NET_201, __A01_NET_202, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1023(__A01_1__F15A, __A01_1__scaler_s15__FS_n, __A01_NET_204, __A01_1__F15B, __A01_NET_203, __A01_1__FS15, GND, __A01_NET_204, __A01_1__FS15, __A01_1__scaler_s15__FS_n, __A01_1__scaler_s15__FS_n, __A01_NET_203, __A01_1__FS15, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1024(__A01_NET_204, __A01_1__F14A, __A01_1__F16A, __A01_1__F15A, __A01_NET_205, __A01_NET_206, GND, __A01_NET_205, __A01_NET_206, __A01_1__F15A, __A01_1__F16B, __A01_NET_203, __A01_1__F15B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1025(__A01_1__F16A, __A01_1__scaler_s16__FS_n, __A01_NET_206, __A01_1__F16B, __A01_NET_205, __A01_1__FS16, GND, __A01_NET_206, __A01_1__FS16, __A01_1__scaler_s16__FS_n, __A01_1__scaler_s16__FS_n, __A01_NET_205, __A01_1__FS16, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1026(F17A, __A01_1__scaler_s17__FS_n, __A01_NET_208, F17B, __A01_NET_207, __A01_1__FS17, GND, __A01_NET_208, __A01_1__FS17, __A01_1__scaler_s17__FS_n, __A01_1__scaler_s17__FS_n, __A01_NET_207, __A01_1__FS17, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1027(F17A, __A01_1__F16A, __A01_NET_208, __A01_1__F16A, F17B, __A01_NET_207, GND,  ,  ,  ,  , __A01_NET_208, __A01_NET_207, VCC, SIM_RST, SIM_CLK);
    U74HC04 U1028(__A01_1__scaler_s2__FS_n, __A01_1__FS02A, __A01_1__scaler_s3__FS_n, __A01_1__FS03A, __A01_1__scaler_s4__FS_n, __A01_1__FS04A, GND, __A01_1__FS05A, __A01_1__scaler_s5__FS_n, F05A_n, __A01_1__F05A, F05B_n, __A01_1__F05B, VCC, SIM_RST, SIM_CLK);
    U74HC02 U1029(__A01_1__CHAT01, RCHAT_n, __A01_1__scaler_s6__FS_n, __A01_1__CHAT02, RCHAT_n, __A01_1__scaler_s7__FS_n, GND, RCHAT_n, __A01_1__scaler_s8__FS_n, __A01_1__CHAT03, RCHAT_n, __A01_1__scaler_s9__FS_n, __A01_1__CHAT04, VCC, SIM_RST, SIM_CLK);
    U74HC02 U1030(__A01_1__CHAT05, RCHAT_n, __A01_1__scaler_s10__FS_n, __A01_1__CHAT06, RCHAT_n, __A01_1__scaler_s11__FS_n, GND, RCHAT_n, __A01_1__scaler_s12__FS_n, __A01_1__CHAT07, RCHAT_n, __A01_1__scaler_s13__FS_n, __A01_1__CHAT08, VCC, SIM_RST, SIM_CLK);
    U74HC02 U1031(__A01_1__CHAT09, RCHAT_n, __A01_1__scaler_s14__FS_n, __A01_1__CHAT10, __A01_NET_143, __A01_1__scaler_s15__FS_n, GND, RCHAT_n, __A01_1__scaler_s16__FS_n, __A01_1__CHAT11, RCHAT_n, __A01_1__scaler_s17__FS_n, __A01_1__CHAT12, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1032(__A01_2__F18A, __A01_2__scaler_s18__FS_n, __A01_NET_210, __A01_2__F18B, __A01_NET_209, __A01_2__FS18, GND, __A01_NET_210, __A01_2__FS18, __A01_2__scaler_s18__FS_n, __A01_2__scaler_s18__FS_n, __A01_NET_209, __A01_2__FS18, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1033(__A01_2__F18A, F17A, __A01_NET_210, F17A, __A01_2__F18B, __A01_NET_209, GND, __A01_NET_212, __A01_2__F19A, __A01_2__F18A, __A01_NET_211, __A01_NET_210, __A01_NET_209, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1034(__A01_2__F19A, __A01_2__scaler_s19__FS_n, __A01_NET_212, __A01_2__F19B, __A01_NET_211, __A01_2__FS19, GND, __A01_NET_212, __A01_2__FS19, __A01_2__scaler_s19__FS_n, __A01_2__scaler_s19__FS_n, __A01_NET_211, __A01_2__FS19, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1035(__A01_NET_212, __A01_2__F18A, __A01_2__F20A, __A01_2__F19A, __A01_NET_213, __A01_NET_214, GND, __A01_NET_213, __A01_NET_214, __A01_2__F19A, __A01_2__F20B, __A01_NET_211, __A01_2__F19B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1036(__A01_2__F20A, __A01_2__scaler_s20__FS_n, __A01_NET_214, __A01_2__F20B, __A01_NET_213, __A01_2__FS20, GND, __A01_NET_214, __A01_2__FS20, __A01_2__scaler_s20__FS_n, __A01_2__scaler_s20__FS_n, __A01_NET_213, __A01_2__FS20, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1037(__A01_2__F21A, __A01_2__scaler_s21__FS_n, __A01_NET_216, __A01_2__F21B, __A01_NET_215, __A01_2__FS21, GND, __A01_NET_216, __A01_2__FS21, __A01_2__scaler_s21__FS_n, __A01_2__scaler_s21__FS_n, __A01_NET_215, __A01_2__FS21, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1038(__A01_2__F21A, __A01_2__F20A, __A01_NET_216, __A01_2__F20A, __A01_2__F21B, __A01_NET_215, GND, __A01_NET_218, __A01_2__F22A, __A01_2__F21A, __A01_NET_217, __A01_NET_216, __A01_NET_215, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1039(__A01_2__F22A, __A01_2__scaler_s22__FS_n, __A01_NET_218, __A01_2__F22B, __A01_NET_217, __A01_2__FS22, GND, __A01_NET_218, __A01_2__FS22, __A01_2__scaler_s22__FS_n, __A01_2__scaler_s22__FS_n, __A01_NET_217, __A01_2__FS22, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1040(__A01_NET_218, __A01_2__F21A, __A01_2__F23A, __A01_2__F22A, __A01_NET_219, __A01_NET_220, GND, __A01_NET_219, __A01_NET_220, __A01_2__F22A, __A01_2__F23B, __A01_NET_217, __A01_2__F22B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1041(__A01_2__F23A, __A01_2__scaler_s23__FS_n, __A01_NET_220, __A01_2__F23B, __A01_NET_219, __A01_2__FS23, GND, __A01_NET_220, __A01_2__FS23, __A01_2__scaler_s23__FS_n, __A01_2__scaler_s23__FS_n, __A01_NET_219, __A01_2__FS23, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1042(__A01_2__F24A, __A01_2__scaler_s24__FS_n, __A01_NET_222, __A01_2__F24B, __A01_NET_221, __A01_2__FS24, GND, __A01_NET_222, __A01_2__FS24, __A01_2__scaler_s24__FS_n, __A01_2__scaler_s24__FS_n, __A01_NET_221, __A01_2__FS24, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1043(__A01_2__F24A, __A01_2__F23A, __A01_NET_222, __A01_2__F23A, __A01_2__F24B, __A01_NET_221, GND, __A01_NET_224, __A01_2__F25A, __A01_2__F24A, __A01_NET_223, __A01_NET_222, __A01_NET_221, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1044(__A01_2__F25A, __A01_2__scaler_s25__FS_n, __A01_NET_224, __A01_2__F25B, __A01_NET_223, __A01_2__FS25, GND, __A01_NET_224, __A01_2__FS25, __A01_2__scaler_s25__FS_n, __A01_2__scaler_s25__FS_n, __A01_NET_223, __A01_2__FS25, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1045(__A01_NET_224, __A01_2__F24A, __A01_2__F26A, __A01_2__F25A, __A01_NET_225, __A01_NET_226, GND, __A01_NET_225, __A01_NET_226, __A01_2__F25A, __A01_2__F26B, __A01_NET_223, __A01_2__F25B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1046(__A01_2__F26A, __A01_2__scaler_s26__FS_n, __A01_NET_226, __A01_2__F26B, __A01_NET_225, __A01_2__FS26, GND, __A01_NET_226, __A01_2__FS26, __A01_2__scaler_s26__FS_n, __A01_2__scaler_s26__FS_n, __A01_NET_225, __A01_2__FS26, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1047(__A01_2__F27A, __A01_2__scaler_s27__FS_n, __A01_NET_228, __A01_2__F27B, __A01_NET_227, __A01_2__FS27, GND, __A01_NET_228, __A01_2__FS27, __A01_2__scaler_s27__FS_n, __A01_2__scaler_s27__FS_n, __A01_NET_227, __A01_2__FS27, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1048(__A01_2__F27A, __A01_2__F26A, __A01_NET_228, __A01_2__F26A, __A01_2__F27B, __A01_NET_227, GND, __A01_NET_230, __A01_2__F28A, __A01_2__F27A, __A01_NET_229, __A01_NET_228, __A01_NET_227, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1049(__A01_2__F28A, __A01_2__scaler_s28__FS_n, __A01_NET_230, __A01_2__F28B, __A01_NET_229, __A01_2__FS28, GND, __A01_NET_230, __A01_2__FS28, __A01_2__scaler_s28__FS_n, __A01_2__scaler_s28__FS_n, __A01_NET_229, __A01_2__FS28, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1050(__A01_NET_230, __A01_2__F27A, __A01_2__F29A, __A01_2__F28A, __A01_NET_231, __A01_NET_232, GND, __A01_NET_231, __A01_NET_232, __A01_2__F28A, __A01_2__F29B, __A01_NET_229, __A01_2__F28B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1051(__A01_2__F29A, __A01_2__scaler_s29__FS_n, __A01_NET_232, __A01_2__F29B, __A01_NET_231, __A01_2__FS29, GND, __A01_NET_232, __A01_2__FS29, __A01_2__scaler_s29__FS_n, __A01_2__scaler_s29__FS_n, __A01_NET_231, __A01_2__FS29, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1052(__A01_2__F30A, __A01_2__scaler_s30__FS_n, __A01_NET_234, __A01_2__F30B, __A01_NET_233, __A01_2__FS30, GND, __A01_NET_234, __A01_2__FS30, __A01_2__scaler_s30__FS_n, __A01_2__scaler_s30__FS_n, __A01_NET_233, __A01_2__FS30, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1053(__A01_2__F30A, __A01_2__F29A, __A01_NET_234, __A01_2__F29A, __A01_2__F30B, __A01_NET_233, GND, __A01_NET_235, __A01_2__F31A, __A01_2__F30A, __A01_NET_236, __A01_NET_234, __A01_NET_233, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1054(__A01_2__F31A, __A01_2__scaler_s31__FS_n, __A01_NET_235, __A01_2__F31B, __A01_NET_236, __A01_2__FS31, GND, __A01_NET_235, __A01_2__FS31, __A01_2__scaler_s31__FS_n, __A01_2__scaler_s31__FS_n, __A01_NET_236, __A01_2__FS31, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1055(__A01_NET_235, __A01_2__F30A, __A01_2__F32A, __A01_2__F31A, __A01_NET_237, __A01_NET_238, GND, __A01_NET_237, __A01_NET_238, __A01_2__F31A, __A01_2__F32B, __A01_NET_236, __A01_2__F31B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1056(__A01_2__F32A, __A01_2__scaler_s32__FS_n, __A01_NET_238, __A01_2__F32B, __A01_NET_237, __A01_2__FS32, GND, __A01_NET_238, __A01_2__FS32, __A01_2__scaler_s32__FS_n, __A01_2__scaler_s32__FS_n, __A01_NET_237, __A01_2__FS32, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U1057(__A01_2__F33A, __A01_2__scaler_s33__FS_n, __A01_NET_240, __A01_2__F33B, __A01_NET_239, __A01_2__FS33, GND, __A01_NET_240, __A01_2__FS33, __A01_2__scaler_s33__FS_n, __A01_2__scaler_s33__FS_n, __A01_NET_239, __A01_2__FS33, VCC, SIM_RST, SIM_CLK);
    U74HC27 U1058(__A01_2__F33A, __A01_2__F32A, __A01_NET_240, __A01_2__F32A, __A01_2__F33B, __A01_NET_239, GND,  ,  ,  ,  , __A01_NET_240, __A01_NET_239, VCC, SIM_RST, SIM_CLK);
    U74HC02 U1059(__A01_2__CHAT13, RCHAT_n, __A01_2__scaler_s18__FS_n, __A01_2__CHAT14, RCHAT_n, __A01_2__scaler_s19__FS_n, GND, RCHBT_n, __A01_2__scaler_s20__FS_n, __A01_2__CHBT01, RCHBT_n, __A01_2__scaler_s21__FS_n, __A01_2__CHBT02, VCC, SIM_RST, SIM_CLK);
    U74HC02 U1060(__A01_2__CHBT03, RCHBT_n, __A01_2__scaler_s22__FS_n, __A01_2__CHBT04, RCHBT_n, __A01_2__scaler_s23__FS_n, GND, RCHBT_n, __A01_2__scaler_s24__FS_n, __A01_2__CHBT05, RCHBT_n, __A01_2__scaler_s25__FS_n, __A01_2__CHBT06, VCC, SIM_RST, SIM_CLK);
    U74HC02 U1061(__A01_2__CHBT07, RCHBT_n, __A01_2__scaler_s26__FS_n, __A01_2__CHBT08, RCHBT_n, __A01_2__scaler_s27__FS_n, GND, RCHBT_n, __A01_2__scaler_s28__FS_n, __A01_2__CHBT09, RCHBT_n, __A01_2__scaler_s29__FS_n, __A01_2__CHBT10, VCC, SIM_RST, SIM_CLK);
    U74HC02 U1062(__A01_2__CHBT11, RCHBT_n, __A01_2__scaler_s30__FS_n, __A01_2__CHBT12, __A01_NET_163, __A01_2__scaler_s31__FS_n, GND, RCHBT_n, __A01_2__scaler_s32__FS_n, __A01_2__CHBT13, RCHBT_n, __A01_2__scaler_s33__FS_n, __A01_2__CHBT14, VCC, SIM_RST, SIM_CLK);
    U74HC04 U1063(F07B, F07B_n, F10A, F10A_n, F09B, F09B_n, GND, FS07_n, __A01_1__FS07, FS07A, FS07_n, FS05_n, __A01_1__FS05, VCC, SIM_RST, SIM_CLK);
    U74HC04 U1064(FS09, FS09_n,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2001(__A02_1__cdiv_1__D, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__B, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__B, __A02_1__cdiv_1__FS, GND, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__A, __A02_1__cdiv_1__FS, __A02_1__cdiv_1__A, __A02_1__cdiv_1__FS, PHS2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U2002(__A02_1__cdiv_1__D, CLOCK, __A02_1__cdiv_1__B, CLOCK, PHS2, __A02_1__cdiv_1__A, GND, __A02_2__EDSET, P02, P03_n, P04, __A02_1__cdiv_1__B, __A02_1__cdiv_1__A, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1) U2003(__A02_1__cdiv_1__D, __A02_1__cdiv_2__F, PHS2, PHS2_n, PHS4, PHS4_n, GND, __A02_NET_127, __A02_1__cdiv_1__B, CT, __A02_NET_127, CT_n, CT, VCC, SIM_RST, SIM_CLK);
    U74HC02 U2004(PHS4, __A02_1__cdiv_2__F, __A02_1__cdiv_1__A, __A02_1__oddset, STOP, __A02_1__RINGA_n, GND, P02_n, P04, __A02_2__SB4, P01, __A02_NET_154, __A02_NET_155, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1) U2005(__A02_1__cdiv_1__FS_n, WT, WT, WT_n, WT, TT_n, GND, __A02_1__ovfstb_r5, __A02_1__ovfstb_r4, __A02_1__ovfstb_r6, __A02_1__ovfstb_r5, __A02_1__OVFSTB_n, __A02_1__ovfstb_r2, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2006(__A02_1__cdiv_2__D, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__FS, GND, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__A, __A02_1__cdiv_2__FS, __A02_1__cdiv_2__A, __A02_1__cdiv_2__FS, __A02_1__cdiv_2__C, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U2007(__A02_1__cdiv_2__D, __A02_1__cdiv_2__F, __A02_1__cdiv_2__B, __A02_1__cdiv_2__F, __A02_1__cdiv_2__C, __A02_1__cdiv_2__A, GND, P03, __A02_2__EDSET, __A02_NET_168, P03_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__A, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U2008(__A02_1__cdiv_2__D, __A02_1__RINGA_n, __A02_1__oddset, __A02_1__ODDSET_n, __A02_1__cdiv_2__C, __A02_1__RINGB_n, GND, __A02_1__evnset, __A02_1__RINGB_n, __A02_1__EVNSET_n, __A02_1__evnset, RT, __A02_1__cdiv_1__A, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U2009(__A02_1__ovfstb_r1, CT_n, __A02_1__ovfstb_r2, __A02_1__ovfstb_r2, __A02_1__ovfstb_r6, __A02_1__ovfstb_r1, GND, __A02_1__ovfstb_r4, __A02_1__ovfstb_r2, __A02_1__ovfstb_r3, __A02_1__ovfstb_r3, __A02_1__ovfstb_r1, __A02_1__ovfstb_r4, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U2010(CT, PHS3_n, WT_n, CLK, WT_n, MONWT, GND, Q2A, WT_n, RT_n, RT, TIMR, __A02_NET_159, VCC, SIM_RST, SIM_CLK);
    U74HC27 U2011(__A02_1__RINGB_n, P05_n, P04, P05, __A02_1__RINGA_n, __A02_NET_166, GND, __A02_NET_148, __A02_2__T12DC_n, __A02_NET_152, __A02_1__EVNSET_n, __A02_NET_164, P04_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2012(P01, __A02_NET_164, P01_n, P01_n, P01, __A02_NET_166, GND, __A02_1__RINGA_n, P01, __A02_NET_169, P01_n, __A02_1__RINGB_n, __A02_NET_167, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2013(P02, __A02_NET_169, P02_n, P02_n, P02, __A02_NET_167, GND, __A02_1__RINGB_n, P02, __A02_NET_168, P02_n, __A02_1__RINGA_n, __A02_NET_162, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2014(__A02_NET_154, __A02_NET_155, STOP_n, P03_n, P03, __A02_NET_162, GND, __A02_1__RINGA_n, P03, __A02_NET_161, P03_n, __A02_1__RINGB_n, __A02_NET_160, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2015(P04, __A02_NET_161, P04_n, P04_n, P04, __A02_NET_160, GND, __A02_1__RINGB_n, P04, __A02_NET_165, P04_n, __A02_1__RINGA_n, __A02_NET_163, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2016(P05, __A02_NET_165, P05_n, P05_n, P05, __A02_NET_163, GND, __A02_NET_152, GOJ1, __A02_NET_153, __A02_1__EVNSET_n, __A02_NET_147, __A02_NET_149, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2017(__A02_2__F01D, FS01_n, __A02_2__F01B, FS01_n, __A02_2__F01B, FS01, GND, FS01_n, __A02_2__F01A, FS01, __A02_2__F01A, FS01, __A02_2__F01C, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U2018(__A02_2__F01D, P01_n, __A02_2__F01B, P01_n, __A02_2__F01C, __A02_2__F01A, GND,  ,  ,  ,  , __A02_2__F01B, __A02_2__F01A, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b1, 1'b0) U2019(SBY, ALGA, STRT1, STRT2, __A02_NET_153, __A02_NET_151, GND, __A02_NET_146, __A02_2__T12DC_n, __A02_NET_141, __A02_1__EVNSET_n, __A02_NET_150, MSTRTP, VCC, SIM_RST, SIM_CLK);
    assign __A02_NET_152 = __A02_NET_152_U2020_2;
    assign __A02_NET_152 = __A02_NET_152_U2020_4;
    U74LVC07 U2020(__A02_NET_150, __A02_NET_152_U2020_2, __A02_NET_151, __A02_NET_152_U2020_4,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0) U2021(__A02_NET_152, __A02_NET_147, MSTP, __A02_NET_141, GOJAM_n, GOJAM, GND, MGOJAM, GOJAM, STOP, STOP_n, MSTPIT_n, STOP, VCC, SIM_RST, SIM_CLK);
    U74HC02 U2022(__A02_NET_142, __A02_1__EVNSET_n, MSTP, GOJAM_n, STRT2, STOPA, GND, STOPA, __A02_NET_144, STOP_n, STRT2, __A02_NET_158, __A02_NET_159, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U2023(__A02_NET_143, __A02_NET_148, STOPA, STOPA, __A02_NET_143, __A02_NET_149, GND, __A02_NET_146, __A02_NET_144, __A02_NET_145, __A02_NET_145, __A02_NET_142, __A02_NET_144, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U2024(__A02_3__T12SET, GOJAM, __A02_3__T01DC_n, __A02_NET_193, GOJAM, __A02_NET_190, GND, __A02_NET_193, __A02_3__T02DC_n, __A02_NET_192, GOJAM, __A02_2__T12DC_n, __A02_NET_191, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U2025(__A02_NET_191, __A02_2__T12DC_n, __A02_NET_190, __A02_NET_181, __A02_2__T12DC_n, __A02_1__ODDSET_n, GND, __A02_2__T12DC_n, __A02_1__EVNSET_n, T12, __A02_NET_181, __A02_NET_190, __A02_3__T01DC_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U2026(__A02_NET_180, __A02_3__T01DC_n, __A02_1__EVNSET_n, T01, __A02_3__T01DC_n, __A02_1__ODDSET_n, GND, __A02_NET_180, __A02_NET_193, __A02_3__T02DC_n, __A02_3__T02DC_n, __A02_1__ODDSET_n, __A02_NET_185, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2027(T02, __A02_3__T02DC_n, __A02_1__EVNSET_n, __A02_3__T03DC_n, __A02_NET_185, __A02_NET_192, GND, __A02_3__T03DC_n, __A02_1__EVNSET_n, __A02_NET_186, __A02_3__T03DC_n, __A02_1__ODDSET_n, T03, VCC, SIM_RST, SIM_CLK);
    U74HC27 U2028(__A02_3__T03DC_n, __A02_NET_188, __A02_3__T04DC_n, __A02_NET_187, GOJAM, __A02_NET_188, GND, __A02_NET_187, __A02_3__T05DC_n, __A02_NET_189, GOJAM, __A02_NET_192, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U2029(__A02_3__T04DC_n, __A02_NET_186, __A02_NET_188, __A02_NET_183, __A02_3__T04DC_n, __A02_1__ODDSET_n, GND, __A02_3__T04DC_n, __A02_1__EVNSET_n, T04, __A02_NET_183, __A02_NET_187, __A02_3__T05DC_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U2030(__A02_NET_174, __A02_3__T05DC_n, __A02_1__EVNSET_n, T05, __A02_3__T05DC_n, __A02_1__ODDSET_n, GND, __A02_NET_189, __A02_NET_174, __A02_3__T06DC_n, __A02_1__EVNSET_n, __A02_3__T06DC_n, T06, VCC, SIM_RST, SIM_CLK);
    U74HC27 U2031(GOJAM, __A02_NET_196, GOJAM, __A02_NET_195, __A02_3__T07DC_n, __A02_NET_196, GND, __A02_NET_195, GOJAM, __A02_NET_198, __A02_3__T08DC_n, __A02_NET_189, __A02_3__T06DC_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2032(__A02_NET_182, __A02_1__ODDSET_n, __A02_3__T06DC_n, __A02_3__T07DC_n, __A02_NET_196, __A02_NET_182, GND, __A02_1__ODDSET_n, __A02_3__T07DC_n, T07, __A02_1__EVNSET_n, __A02_3__T07DC_n, __A02_NET_184, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U2033(__A02_3__T08DC_n, __A02_NET_195, __A02_NET_184, T08, __A02_1__EVNSET_n, __A02_3__T08DC_n, GND, __A02_1__ODDSET_n, __A02_3__T08DC_n, __A02_NET_176, __A02_NET_198, __A02_NET_176, __A02_3__T09DC_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U2034(GOJAM, __A02_NET_197, GOJAM, __A02_NET_194, __A02_3__T10DC_n, __A02_NET_197, GND, __A02_NET_194, GOJAM, __A02_NET_177, __A02_NET_179, __A02_NET_198, __A02_3__T09DC_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U2035(T09, __A02_1__ODDSET_n, __A02_3__T09DC_n, __A02_NET_175, __A02_1__EVNSET_n, __A02_3__T09DC_n, GND, __A02_NET_197, __A02_NET_175, __A02_3__T10DC_n, __A02_1__EVNSET_n, __A02_NET_197, __A02_NET_177, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2036(__A02_NET_178, __A02_1__ODDSET_n, __A02_3__T10DC_n, __A02_NET_179, __A02_NET_194, __A02_NET_178, GND, __A02_1__EVNSET_n, __A02_3__T10DC_n, T10, __A02_1__ODDSET_n, __A02_NET_179, T11, VCC, SIM_RST, SIM_CLK);
    U74HC02 U2037(__A02_NET_170, __A02_NET_193, __A02_NET_190, __A02_2__SB0, P02_n, P05, GND, P05_n, P03_n, __A02_2__SB1, P05_n, P02, SB2, VCC, SIM_RST, SIM_CLK);
    U74HC27 U2038(__A02_NET_187, __A02_NET_188, __A02_NET_198, __A02_NET_197, __A02_1__EVNSET_n, __A02_NET_172, GND, __A02_NET_173, __A02_NET_189, __A02_NET_196, __A02_NET_195, __A02_NET_171, __A02_NET_192, VCC, SIM_RST, SIM_CLK);
    assign __A02_3__T12SET = __A02_3__T12SET_U2039_2;
    assign __A02_3__T12SET = __A02_3__T12SET_U2039_4;
    assign __A02_3__T12SET = __A02_3__T12SET_U2039_6;
    assign __A02_3__T12SET = __A02_3__T12SET_U2039_8;
    U74LVC07 U2039(__A02_NET_170, __A02_3__T12SET_U2039_2, __A02_NET_171, __A02_3__T12SET_U2039_4, __A02_NET_172, __A02_3__T12SET_U2039_6, GND, __A02_3__T12SET_U2039_8, __A02_NET_173,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0) U2040(T01, T01_n, T01_n, MT01, T02, T02_n, GND, MT02, T02_n, T03_n, T03, MT03, T03_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0) U2041(T04, T04_n, T04_n, MT04, T05, T05_n, GND, MT05, T05_n, T06_n, T06, MT06, T06_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0) U2042(T07, T07_n, T07_n, MT07, T08, T08_n, GND, MT08, T08_n, T09_n, T09, MT09, T09_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0) U2043(T10, T10_n, T10_n, MT10, T11, T11_n, GND, MT11, T11_n, T12_n, T12, MT12, T12_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U2044(WL15_n, WL16, __A02_1__OVFSTB_n, WL15, WL16_n, __A02_3__UNF, GND,  ,  ,  ,  , __A02_3__OVF, __A02_1__OVFSTB_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0) U2045(__A02_3__OVF, OVF_n, __A02_3__UNF, UNF_n, __A02_2__SB0, SB0_n, GND, SB1_n, __A02_2__SB1, SB2_n, SB2, T12A, T12_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U2046(__A02_NET_158, P04, P05_n, __A02_NET_155, STOP_n,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U3001(__A03_NET_166, NISQ, __A03_1__NISQL, __A03_NET_167, STRTFC, __A03_NET_168, GND, RT_n, __A03_NET_163, RBSQ, __A03_NET_163, WT_n, __A03_1__wsqg, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3002(__A03_NET_166, __A03_1__INKBT1, T12_n, __A03_NET_166, __A03_1__RPTFRC, __A03_NET_168, GND, __A03_1__CSQG, T12_n, CT_n, __A03_NET_167, __A03_1__NISQL, STRTFC, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1) U3003(__A03_1__NISQL, NISQL_n, __A03_NET_168, __A03_NET_163, __A03_1__wsqg, __A03_1__WSQG_n, GND, STRTFC, __A03_NET_161, SQEXT, __A03_NET_175, SQEXT_n, __A03_NET_174, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3004(__A03_NET_197, WL16_n, __A03_1__WSQG_n, __A03_NET_210, WL14_n, __A03_1__WSQG_n, GND, WL13_n, __A03_1__WSQG_n, __A03_NET_209,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U3005(__A03_NET_161, GOJAM, MTCSAI, __A03_NET_165, NISQL_n, T12_n, GND, STRTFC, __A03_NET_165, __A03_NET_172, __A03_NET_172, __A03_NET_164, __A03_NET_171, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U3006(EXTPLS, EXT, __A03_NET_164, __A03_1__INKBT1, STRTFC, FUTEXT, GND, __A03_NET_175, __A03_1__RPTFRC, __A03_NET_171, __A03_NET_174, __A03_NET_164, FUTEXT, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b1) U3007(__A03_NET_170, __A03_NET_172, FUTEXT, __A03_NET_174, __A03_NET_175, __A03_NET_170, GND, INHPLS, __A03_1__INHINT, __A03_NET_169, KRPT, IIP, IIP_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U3008(__A03_NET_175, __A03_1__MSQEXT, __A03_NET_169, __A03_1__MINHL, IIP_n, __A03_1__MIIP, GND, __A03_1__MSQ16, __A03_NET_202, __A03_1__MSQ14, __A03_NET_188, __A03_1__MSQ13, __A03_NET_190, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3009(__A03_NET_169, RELPLS, IIP_n, GOJAM, n5XP4, IIP, GND, __A03_NET_196, FUTEXT, NISQL_n, T12_n, __A03_1__INHINT, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3010(PHS2_n, RUPTOR_n, OVNHRP, __A03_1__INHINT, IIP, __A03_NET_194, GND, __A03_NET_192, __A03_NET_193, STRTFC, T02, __A03_NET_195, MNHRPT, VCC, SIM_RST, SIM_CLK);
    assign RPTSET = RPTSET_U3011_2;
    assign RPTSET = RPTSET_U3011_4;
    assign RPTSET = RPTSET_U3011_6;
    U74LVC07 U3011(__A03_NET_196, RPTSET_U3011_2, __A03_NET_195, RPTSET_U3011_4, __A03_NET_194, RPTSET_U3011_6, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b1) U3012(__A03_NET_193, RPTSET, __A03_NET_192, __A03_NET_202, __A03_NET_197, __A03_1__SQR16, GND, __A03_NET_210, __A03_1__SQR14, __A03_NET_188, __A03_NET_209, __A03_1__SQR13, __A03_NET_190, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3013(__A03_NET_202, __A03_1__RPTFRC, __A03_NET_188, __A03_1__RPTFRC, __A03_1__CSQG, __A03_1__SQR14, GND, __A03_1__SQR13, __A03_NET_190, __A03_1__RPTFRC, __A03_1__CSQG, __A03_1__SQR16, __A03_1__CSQG, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U3014(__A03_NET_200, __A03_NET_202, INKL, __A03_NET_199, INKL, __A03_1__SQR16, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U3015(__A03_NET_189, __A03_NET_187, __A03_NET_190, __A03_NET_187, __A03_NET_203, __A03_NET_201, GND, __A03_NET_208, __A03_NET_189, __A03_NET_188, __A03_NET_203, __A03_NET_198, __A03_NET_203, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3016(__A03_NET_190, __A03_NET_188, __A03_NET_189, __A03_NET_187, __A03_NET_186, __A03_NET_206, GND, __A03_NET_178, __A03_NET_190, __A03_NET_187, __A03_NET_186, __A03_NET_207, __A03_NET_203, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U3017(__A03_NET_189, __A03_NET_186, __A03_NET_190, __A03_NET_188, __A03_NET_186, __A03_NET_204, GND, __A03_NET_191, __A03_1__RPTFRC, __A03_NET_185, __A03_1__SQR12, __A03_NET_205, __A03_NET_188, VCC, SIM_RST, SIM_CLK);
    U74HC04 U3018(__A03_NET_201, SQ1_n, __A03_NET_208, SQ2_n, __A03_NET_207, __A03_1__SQ3_n, GND, __A03_1__SQ4_n, __A03_NET_206, __A03_1__SQ6_n, __A03_NET_205, __A03_1__SQ7_n, __A03_NET_204, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3019(__A03_NET_185, WL12_n, __A03_1__WSQG_n, __A03_NET_177, WL11_n, __A03_1__WSQG_n, GND, __A03_NET_191, __A03_1__CSQG, __A03_1__SQR12, __A03_NET_176, __A03_1__CSQG, __A03_1__SQR11, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b1, 1'b0) U3020(__A03_1__RPTFRC, __A03_NET_177, __A03_1__RPTFRC, __A03_NET_184, __A03_NET_183, __A03_NET_182, GND, __A03_1__INKBT1, INKL, T01_n, STD2, __A03_NET_176, __A03_1__SQR11, VCC, SIM_RST, SIM_CLK);
    U74HC04 U3021(__A03_NET_191, __A03_1__MSQ12, __A03_NET_176, __A03_1__MSQ11, __A03_NET_182, __A03_1__MSQ10, GND, SQR12_n, __A03_1__SQR12, __A03_1__RPTFRC, __A03_NET_193, __A03_1__SQ5_n, __A03_NET_178, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3022(__A03_1__QC0, __A03_1__SQR11, __A03_1__SQR12, __A03_NET_181, __A03_NET_176, __A03_1__SQR12, GND, __A03_1__SQR11, __A03_NET_191, __A03_NET_180, __A03_NET_191, __A03_NET_176, __A03_NET_179, VCC, SIM_RST, SIM_CLK);
    U74HC04 U3023(__A03_1__QC0, QC0_n, __A03_NET_181, QC1_n, __A03_NET_180, QC2_n, GND, QC3_n, __A03_NET_179, SQR10, __A03_NET_182, SQR10_n, __A03_NET_183, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3024(__A03_NET_184, WL10_n, __A03_1__WSQG_n, __A03_NET_183, __A03_NET_182, __A03_1__CSQG, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U3025(__A03_NET_200, __A03_NET_186, __A03_NET_199, __A03_NET_203, __A03_NET_188, __A03_NET_187, GND, __A03_NET_189, __A03_NET_190, SQ0_n, __A03_NET_198, MP3A, MP3_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3026(__A03_NET_225, __A03_1__SQ5_n, QC0_n, __A03_NET_226, __A03_1__SQ5_n, SQEXT_n, GND, __A03_NET_225, __A03_NET_226, __A03_NET_227, __A03_NET_227, ST0_n, IC1, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1) U3027(__A03_NET_225, __A03_2__SQ5QC0_n, IC2, IC2_n, __A03_NET_233, EXST1_n, GND, TC0_n, TC0, IC3, __A03_2__IC3_n, __A03_2__NEXST0_n, __A03_2__NEXST0, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3028(IC2, __A03_NET_227, ST1_n, __A03_NET_229, SQEXT_n, __A03_1__QC0, GND, SQEXT_n, ST1_n, __A03_NET_233, __A03_NET_233, __A03_2__NEXST0, __A03_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3029(__A03_NET_229, __A03_1__SQ6_n, SQ1_n, __A03_2__NEXST0_n, __A03_1__QC0, TCF0, GND, __A03_2__IC3_n, TC0, STD2, TCF0, IC11, ST0_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3030(IC6, __A03_NET_232, __A03_1__SQ3_n, IC7, __A03_NET_232, __A03_1__SQ4_n, GND, SQ0_n, __A03_2__NEXST0_n, TC0, SQEXT, ST0_n, __A03_2__NEXST0, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3031(DCS0, __A03_1__SQ4_n, EXST0_n, DCA0, EXST0_n, __A03_1__SQ3_n, GND, DCS0, DCA0, __A03_2__IC4_n, QC1_n, ST1_n, __A03_NET_216, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3032(IC7, IC6, IC1, DCS0, DCA0, __A03_NET_221, GND, IC5, __A03_NET_214, __A03_1__SQ5_n, SQEXT, __A03_NET_220, IC11, VCC, SIM_RST, SIM_CLK);
    assign __A03_2__IC13_n = __A03_2__IC13_n_U3033_2;
    assign __A03_2__IC13_n = __A03_2__IC13_n_U3033_4;
    U74LVC07 U3033(__A03_NET_220, __A03_2__IC13_n_U3033_2, __A03_NET_221, __A03_2__IC13_n_U3033_4,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U3034(__A03_2__IC4_n, IC4, __A03_2__IC13_n, IC13, IC5, IC5_n, GND, IC9, __A03_2__IC9_n, QXCH0_n, __A03_2__QXCH0, EXST0_n, __A03_NET_213, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3035(__A03_NET_215, QC3_n, ST0_n, __A03_NET_214, __A03_NET_216, __A03_NET_215, GND, __A03_2__LXCH0, DXCH0, IC8_n, ST0_n, SQEXT_n, __A03_NET_213, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3036(__A03_2__NEXST0_n, QC1_n, SQ2_n, QC1_n, EXST0_n, __A03_2__QXCH0, GND, TS0, __A03_1__SQ5_n, QC2_n, __A03_2__NEXST0_n, __A03_2__LXCH0, SQ2_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U3037(__A03_2__IC9_n, IC5, TS0, __A03_2__QXCH0, __A03_2__LXCH0,  , GND,  , SQ2_n, QC0_n, SQEXT, ST1_n, __A03_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC04 U3038(TS0, TS0_n, IC10_n, IC10, DAS0, DAS0_n, GND, __A03_2__BZF0_n, __A03_2__BZF0, __A03_2__BMF0_n, __A03_2__BMF0, IC16, IC16_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3039(__A03_1__SQ5_n, __A03_2__NEXST0_n, SQ2_n, __A03_2__NEXST0_n, QC0_n, DAS0, GND, IC10_n, IC4, DXCH0, DAS0, DXCH0, QC1_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3040(SQ1_n, __A03_1__QC0, EXST0_n, __A03_1__QC0, __A03_1__SQ6_n, __A03_2__BMF0, GND, CCS0, SQ1_n, QC0_n, __A03_2__NEXST0_n, __A03_2__BZF0, EXST0_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3041(IC15_n, __A03_2__BMF0, __A03_2__BZF0, __A03_NET_217, __A03_2__BZF0_n, BR2_n, GND, __A03_2__BMF0_n, BR1B2B, __A03_NET_218, __A03_NET_217, __A03_NET_218, IC16_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U3042(IC17, IC16, IC15_n, DAS1_n, __A03_NET_212, ADS0, GND, CCS0, MSU0, IC12_n, __A03_1__SQ7_n, __A03_2__NEXST0_n, MASK0, VCC, SIM_RST, SIM_CLK);
    U74HC04 U3043(IC15_n, IC15, CCS0, CCS0_n, DAS1_n, DAS1, GND, IC12, IC12_n, MSU0_n, MSU0, AUG0_n, __A03_2__AUG0, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U3044(SQ2_n, QC3_n, QC2_n, SQ2_n, __A03_2__NEXST0_n, INCR0, GND, MSU0, SQ2_n, EXST0_n, QC0_n, ADS0, __A03_2__NEXST0_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3045(SQ2_n, EXST0_n, SQ2_n, EXST0_n, QC3_n, __A03_2__DIM0, GND, MP3, ST3_n, __A03_1__SQ7_n, SQEXT_n, __A03_2__AUG0, QC2_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U3046(__A03_2__DIM0, DIM0_n, MP3, MP3_n, MP1, MP1_n, GND, MP0_n, MP0, TCSAJ3_n, TCSAJ3, RSM3_n, RSM3, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3047(ST1_n, __A03_1__SQ7_n, ST0_n, __A03_1__SQ7_n, SQEXT_n, MP0, GND, TCSAJ3, SQ0_n, SQEXT, ST3_n, MP1, SQEXT_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U3048(ST3_n, __A03_2__SQ5QC0_n, __A03_1__SQ6_n, EXST0_n, QC0_n, SU0, GND, __A03_NET_219, MP0, MASK0, RXOR0, RSM3, SQEXT, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0) U3049(MASK0, MASK0_n, __A03_NET_219, IC14, __A03_2__NDX0, NDX0_n, GND, NDXX1_n, __A03_2__NDXX1, GOJ1_n, GOJ1, IC11_n, IC11, VCC, SIM_RST, SIM_CLK);
    U74HC02 U3050(AD0, __A03_2__NEXST0_n, __A03_1__SQ6_n,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U3051(__A03_2__NEXST0_n, __A03_1__SQ5_n, SQEXT_n, __A03_1__SQ5_n, ST1_n, __A03_2__NDXX1, GND, GOJ1, SQEXT, ST1_n, SQ0_n, __A03_2__NDX0, QC0_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U4001(T12USE_n, DVST, __A04_NET_243, DIVSTG, T12USE_n, T03_n, GND, __A04_NET_244, __A04_NET_242, __A04_NET_268, GOJAM, MTCSAI, __A04_NET_249, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U4002(T03_n, T12USE_n, T12USE_n, RSTSTG, GOJAM, __A04_NET_243, GND, __A04_NET_242, PHS3_n, __A04_NET_243, T12_n, __A04_NET_244, PHS3_n, VCC, SIM_RST, SIM_CLK);
    assign __A04_NET_250 = __A04_NET_250_U4003_2;
    assign __A04_NET_250 = __A04_NET_250_U4003_4;
    assign __A04_NET_238 = __A04_NET_238_U4003_6;
    assign __A04_NET_238 = __A04_NET_238_U4003_8;
    assign __A04_1__SGUM = __A04_1__SGUM_U4003_10;
    assign __A04_1__SGUM = __A04_1__SGUM_U4003_12;
    U74LVC07 U4003(__A04_NET_249, __A04_NET_250_U4003_2, __A04_NET_248, __A04_NET_250_U4003_4, __A04_NET_229, __A04_NET_238_U4003_6, GND, __A04_NET_238_U4003_8, __A04_NET_232, __A04_1__SGUM_U4003_10, __A04_NET_198, __A04_1__SGUM_U4003_12, __A04_NET_197, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b1, 1'b0) U4004(ST1, __A04_NET_245, __A04_1__STG1, __A04_1__STG3, __A04_1__STG2, __A04_NET_231, GND, __A04_NET_254, __A04_1__STG2, __A04_1__STG3, __A04_NET_236, __A04_NET_248, __A04_NET_247, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4005(__A04_NET_247, __A04_NET_250, T01, __A04_NET_245, __A04_NET_234, __A04_1__STG3, GND, __A04_NET_268, __A04_NET_250, __A04_NET_241, __A04_NET_247, __A04_NET_268, __A04_NET_246, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U4006(__A04_NET_236, __A04_NET_241, __A04_1__STG1, __A04_1__STG1, __A04_NET_236, __A04_NET_246, GND, ST2, __A04_NET_230, __A04_NET_229, __A04_NET_234, __A04_NET_236, __A04_NET_235, VCC, SIM_RST, SIM_CLK);
    U74HC04 U4007(__A04_NET_236, __A04_1__MST1, __A04_NET_259, __A04_1__MST2, __A04_NET_269, __A04_1__MST3, GND, __A04_1__MBR1, __A04_NET_216, __A04_1__MBR2, __A04_NET_212, __A04_NET_234, DVST, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0) U4008(__A04_NET_231, ST0_n, __A04_NET_254, ST1_n, __A04_NET_264, ST3_n, GND, __A04_1__ST4_n, __A04_NET_252, __A04_1__ST376_n, __A04_1__ST376, DV1376_n, DV1376, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U4009(__A04_NET_235, MTCSAI, __A04_NET_238, GOJAM, T01, __A04_NET_233, GND, __A04_NET_264, __A04_1__STG3, __A04_NET_259, __A04_NET_236, __A04_NET_232, __A04_NET_233, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U4010(__A04_NET_230, __A04_NET_209, XT1_n, XB7_n, NDR100_n,  , GND,  , __A04_NET_256, STRTFC, T01, RSTSTG, __A04_NET_261, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U4011(__A04_NET_262, __A04_NET_268, __A04_NET_238, __A04_NET_237, __A04_NET_233, __A04_NET_268, GND, __A04_NET_262, __A04_1__STG2, __A04_NET_259, __A04_NET_259, __A04_NET_237, __A04_1__STG2, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U4012(__A04_NET_260, __A04_NET_234, __A04_NET_259, __A04_NET_256, __A04_NET_260, __A04_NET_261, GND, __A04_NET_268, __A04_NET_256, __A04_NET_265, __A04_NET_261, __A04_NET_268, __A04_NET_266, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U4013(__A04_NET_269, __A04_NET_265, __A04_1__STG3, __A04_1__STG3, __A04_NET_269, __A04_NET_266, GND, __A04_1__STG1, __A04_1__STG3, __A04_NET_251, __A04_NET_259, __A04_NET_251, __A04_1__ST376, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U4014(STD2, INKL, __A04_1__STG1, __A04_1__STG3, __A04_NET_259,  , GND,  , SQ0_n, EXST1_n, QC3_n, SQR10_n, RUPT1, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4015(__A04_NET_269, __A04_1__STG1, QC0_n, SQEXT_n, SQ1_n, __A04_NET_253, GND, __A04_NET_198, SUMB16_n, SUMA16_n, TSGU_n, __A04_NET_252, __A04_1__STG2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4016(__A04_NET_255, __A04_NET_252, __A04_1__ST376, DV3764, DIV_n, __A04_NET_255, GND, __A04_NET_254, __A04_1__ST376, __A04_1__ST1376_n, DIV_n, __A04_1__ST1376_n, DV1376, VCC, SIM_RST, SIM_CLK);
    U74HC04 U4017(__A04_NET_253, DIV_n, __A04_1__DV0, __A04_1__DV0_n, DV1, DV1_n, GND, DV376_n, __A04_1__DV376, __A04_NET_189, TL15, BR1, __A04_NET_216, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4018(__A04_1__DV0, DIV_n, ST0_n, DV1, DIV_n, ST1_n, GND, DIV_n, __A04_1__ST4_n, DV4, DIV_n, __A04_1__ST376_n, __A04_1__DV376, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4019(__A04_NET_185, SUMA16_n, SUMB16_n, __A04_NET_197, PHS4, PHS3_n, GND, UNF_n, TOV_n, __A04_NET_187, L15_n, __A04_NET_189, __A04_NET_193, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U4020(PHS4_n, WL16_n, __A04_NET_193, __A04_NET_188, __A04_NET_217, __A04_NET_195, GND, __A04_NET_194, __A04_NET_216, __A04_NET_192, __A04_NET_191, __A04_NET_188, TSGN_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4021(__A04_NET_192, TSGN_n, PHS3_n, __A04_NET_191, __A04_NET_189, PHS3_n, GND, TOV_n, PHS2_n, __A04_NET_204, __A04_1__SGUM, __A04_NET_187, __A04_NET_186, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U4022(__A04_NET_196, __A04_NET_185, PHS3_n, TSGU_n, PHS4,  , GND,  , WL16_n, WL15_n, WL14_n, WL13_n, __A04_NET_213, VCC, SIM_RST, SIM_CLK);
    assign __A04_NET_216 = __A04_NET_216_U4023_2;
    assign __A04_NET_216 = __A04_NET_216_U4023_4;
    assign __A04_NET_217 = __A04_NET_217_U4023_6;
    assign __A04_NET_217 = __A04_NET_217_U4023_8;
    assign __A04_NET_222 = __A04_NET_222_U4023_10;
    assign __A04_NET_222 = __A04_NET_222_U4023_12;
    U74LVC07 U4023(__A04_NET_186, __A04_NET_216_U4023_2, __A04_NET_195, __A04_NET_216_U4023_4, __A04_NET_194, __A04_NET_217_U4023_6, GND, __A04_NET_217_U4023_8, __A04_NET_190, __A04_NET_222_U4023_10, __A04_NET_213, __A04_NET_222_U4023_12, __A04_NET_221, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U4024(__A04_NET_190, __A04_NET_204, __A04_NET_196, __A04_NET_201, TOV_n, OVF_n, GND, __A04_NET_208, PHS3_n, __A04_NET_205, TMZ_n, PHS4_n, __A04_NET_220, VCC, SIM_RST, SIM_CLK);
    U74HC04 U4025(__A04_NET_217, BR1_n, __A04_1__TSGN2, __A04_NET_208, __A04_NET_212, BR2, GND, BR2_n, __A04_NET_202, DV4_n, DV4, __A04_NET_332, __A04_NET_331, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4026(GEQZRO_n, PHS4_n, WL16_n, PHS4_n, __A04_NET_208, __A04_NET_210, GND, __A04_NET_203, __A04_NET_210, __A04_NET_222, __A04_NET_202, __A04_NET_199, TPZG_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U4027(__A04_NET_221, WL12_n, WL11_n, WL10_n, WL09_n,  , GND,  , WL08_n, WL07_n, WL06_n, WL05_n, __A04_NET_218, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b0, 1'b1) U4028(__A04_NET_219, WL04_n, WL03_n, WL02_n, WL01_n,  , GND,  , __A04_NET_212, __A04_NET_205, __A04_NET_211, __A04_NET_204, __A04_NET_202, VCC, SIM_RST, SIM_CLK);
    assign __A04_NET_222 = __A04_NET_222_U4029_2;
    assign __A04_NET_222 = __A04_NET_222_U4029_4;
    assign __A04_NET_222 = __A04_NET_222_U4029_6;
    assign __A04_NET_212 = __A04_NET_212_U4029_8;
    assign __A04_NET_212 = __A04_NET_212_U4029_10;
    U74LVC07 U4029(__A04_NET_218, __A04_NET_222_U4029_2, __A04_NET_219, __A04_NET_222_U4029_4, __A04_NET_220, __A04_NET_222_U4029_6, GND, __A04_NET_212_U4029_8, __A04_NET_200, __A04_NET_212_U4029_10, __A04_NET_203,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U4030(__A04_NET_211, TMZ_n, PHS3_n, __A04_NET_200, __A04_NET_199, __A04_NET_201, GND, SQ0_n, EXST0_n, __A04_NET_331, QC3_n, SQEXT, __A04_NET_278, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4031(__A04_NET_332, SQR10, QC0_n, __A04_NET_332, SQR10_n, __A04_2__WRITE0, GND, RAND0, SQR10, __A04_NET_332, QC1_n, READ0, QC0_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U4032(READ0, __A04_2__READ0_n, __A04_2__WRITE0, __A04_2__WRITE0_n, WOR0, __A04_2__WOR0_n, GND, RXOR0_n, RXOR0, __A04_2__RUPT0_n, RUPT0, __A04_2__RUPT1_n, RUPT1, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4033(QC1_n, SQR10_n, SQR10, __A04_NET_332, QC2_n, ROR0, GND, WOR0, QC2_n, __A04_NET_332, SQR10_n, WAND0, __A04_NET_332, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4034(SQR10, __A04_NET_332, QC3_n, __A04_NET_332, SQR10_n, RUPT0, GND, __A04_NET_276, ST0_n, SQR12_n, SQ2_n, RXOR0, QC3_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U4035(__A04_NET_276, __A04_NET_277, INOUT, INOUT_n, __A04_NET_283, __A04_NET_317, GND, BR1B2_n, __A04_2__BR1B2, BR12B_n, __A04_2__BR12B, BR1B2B_n, BR1B2B, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4036(PRINC, __A04_NET_278, __A04_NET_277, RRPA, T03_n, __A04_2__RUPT1_n, GND, T03_n, RXOR0_n, n3XP7, __A04_NET_272, T03_n, __A04_NET_275, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4037(EXST0_n, SQ0_n, INOUT, DV4, PRINC, __A04_NET_312, GND, __A04_NET_327, __A04_NET_275, __A04_NET_273, __A04_NET_280, INOUT, RUPT0, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4038(__A04_NET_272, ROR0, WOR0, __A04_NET_274, T03_n, __A04_NET_271, GND, RAND0, WAND0, __A04_NET_271, DV4_n, T05_n, n5XP28, VCC, SIM_RST, SIM_CLK);
    assign RB_n = RB_n_U4039_2;
    assign RC_n = RC_n_U4039_4;
    assign n5XP11 = n5XP11_U4039_6;
    assign n5XP11 = n5XP11_U4039_8;
    assign RA_n = RA_n_U4039_10;
    assign WG_n = WG_n_U4039_12;
    U74LVC07 U4039(__A04_NET_327, RB_n_U4039_2, __A04_NET_326, RC_n_U4039_4, __A04_NET_329, n5XP11_U4039_6, GND, n5XP11_U4039_8, __A04_NET_328, RA_n_U4039_10, __A04_NET_330, WG_n_U4039_12, __A04_NET_300, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U4040(__A04_NET_274, __A04_NET_285, T05_n, INOUT_n, READ0, __A04_NET_329, GND, WCH_n, __A04_NET_286, n7XP14, __A04_NET_284, __A04_NET_326, __A04_NET_282, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4041(__A04_NET_328, __A04_2__WRITE0, RXOR0, __A04_NET_273, __A04_2__READ0_n, T05_n, GND, __A04_2__WRITE0_n, T05_n, __A04_NET_286, T05_n, __A04_2__WOR0_n, __A04_NET_284, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4042(__A04_NET_285, T05_n, RXOR0_n, __A04_NET_281, T02_n, __A04_2__WRITE0_n, GND, T02_n, INOUT_n, n2XP3, T09_n, __A04_2__RUPT0_n, n9XP1, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4043(__A04_NET_286, __A04_NET_285, RUPT1, IC13, IC12, __A04_NET_287, GND, __A04_NET_300, n9XP1, __A04_NET_282, __A04_NET_280, __A04_NET_330, n2XP3, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4044(__A04_NET_282, T09_n, RXOR0_n, __A04_NET_280, T09_n, __A04_NET_287, GND, __A04_NET_285, __A04_NET_281, __A04_NET_337, T01_n, __A04_2__RUPT1_n, RB2, VCC, SIM_RST, SIM_CLK);
    assign WG_n = WG_n_U4045_2;
    assign __A04_NET_283 = __A04_NET_283_U4045_4;
    assign __A04_NET_283 = __A04_NET_283_U4045_6;
    assign RA_n = RA_n_U4045_8;
    assign WG_n = WG_n_U4045_10;
    assign TMZ_n = TMZ_n_U4045_12;
    U74LVC07 U4045(__A04_NET_337, WG_n_U4045_2, __A04_NET_335, __A04_NET_283_U4045_4, __A04_NET_336, __A04_NET_283_U4045_6, GND, RA_n_U4045_8, __A04_NET_314, WG_n_U4045_10, __A04_NET_302, TMZ_n_U4045_12, __A04_NET_322, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4046(RUPT0, RUPT1, INOUT, MP1, MP3A, __A04_NET_335, GND, __A04_NET_336, __A04_1__DV0, IC15, DV1376, __A04_NET_279, RSM3, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4047(R15, __A04_NET_279, T01_n, n1XP10, T01_n, __A04_1__DV0_n, GND, MP0_n, T03_n, __A04_NET_270, INOUT_n, T03_n, __A04_NET_320, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4048(T02_n, __A04_1__DV0_n, BRDIF_n, TS0_n, T04_n, __A04_NET_299, GND, __A04_NET_294, T04_n, BR1, MP0_n, n2XP5, BR1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4049(n3XP2, T03_n, TS0_n, __A04_2__BR1B2, BR1, BR2_n, GND, BR1_n, BR2, __A04_2__BR12B, __A04_2__BR1B2, __A04_2__BR12B, BRDIF_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4050(BR1B2B, BR2, BR1, n4XP5, TS0_n, T04_n, GND, T04_n, INOUT_n, n4XP11, T04_n, MP3_n, __A04_NET_323, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4051(MP0_n, BR1_n, DV1_n, T04_n, BR2_n, __A04_NET_289, GND, __A04_NET_292, TS0_n, T05_n, BR1B2_n, __A04_NET_319, T04_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4052(T05_n, TS0_n, T07_n, BR1_n, MP3_n, n7XP19, GND, n8XP6, T08_n, DV1_n, BR2, __A04_NET_311, BR12B_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4053(B15X, T05_n, DV1_n, n5XP4, T05_n, RSM3_n, GND, T06_n, DV1_n, n6XP5, T06_n, MP3_n, TL15, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4054(__A04_1__TSGN2, T07_n, MP0_n, __A04_NET_308, T07_n, DV1_n, GND, T08_n, DV1_n, n8XP5, T09_n, MP3_n, __A04_NET_313, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4055(T09_n, BR1, T09_n, MP0_n, BR1_n, __A04_NET_295, GND, __A04_NET_298, MP0_n, T09_n, BRDIF_n, __A04_NET_318, MP0_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4056(KRPT, T09_n, __A04_2__RUPT1_n, MP0T10, T10_n, MP0_n, GND, __A04_NET_317, T02_n, __A04_NET_315, STORE1_n, T09_n, __A04_NET_303, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4057(BR1_n, MP0_n, n1XP10, n8XP5, __A04_NET_313, __A04_NET_314, GND,  ,  ,  ,  , __A04_NET_316, T11_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0) U4058(RSC_n, __A04_2__MRSC, __A04_NET_316, __A04_NET_310, TRSM, __A04_NET_209, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b1) U4059( ,  , __A04_NET_320, B15X, n7XP19, __A04_NET_325, GND, __A04_NET_324, n8XP5, __A04_NET_318, __A04_NET_295,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U4060(__A04_NET_322, n2XP5, n1XP10, __A04_NET_297, __A04_NET_299, __A04_NET_298, GND, n1XP10, MP0T10, __A04_NET_290, __A04_NET_292, __A04_NET_316, __A04_NET_291, VCC, SIM_RST, SIM_CLK);
    assign WY_n = WY_n_U4061_2;
    assign WY_n = WY_n_U4061_4;
    assign WL_n = WL_n_U4061_6;
    assign RC_n = RC_n_U4061_8;
    assign RB_n = RB_n_U4061_10;
    assign CI_n = CI_n_U4061_12;
    U74LVC07 U4061(__A04_NET_325, WY_n_U4061_2, __A04_NET_324, WY_n_U4061_4, __A04_NET_321, WL_n_U4061_6, GND, RC_n_U4061_8, __A04_NET_296, RB_n_U4061_10, __A04_NET_293, CI_n_U4061_12, __A04_NET_297, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U4062(__A04_NET_294, __A04_NET_319, __A04_NET_319, n2XP5, __A04_NET_295, __A04_NET_296, GND, __A04_NET_293, __A04_NET_294, n7XP19, __A04_NET_318, __A04_NET_321, n6XP5, VCC, SIM_RST, SIM_CLK);
    assign TSGN_n = TSGN_n_U4063_2;
    assign TSGN_n = TSGN_n_U4063_4;
    assign RB1_n = RB1_n_U4063_6;
    assign L16_n = L16_n_U4063_8;
    assign R1C_n = R1C_n_U4063_10;
    assign n8PP4 = n8PP4_U4063_12;
    U74LVC07 U4063(__A04_NET_290, TSGN_n_U4063_2, __A04_NET_288, TSGN_n_U4063_4, __A04_NET_291, RB1_n_U4063_6, GND, L16_n_U4063_8, __A04_NET_310, R1C_n_U4063_10, __A04_NET_309, n8PP4_U4063_12, __A04_NET_312, VCC, SIM_RST, SIM_CLK);
    U74HC27 U4064(__A04_NET_289, __A04_NET_270,  ,  ,  ,  , GND,  ,  ,  ,  , __A04_NET_288, __A04_NET_308, VCC, SIM_RST, SIM_CLK);
    U74HC02 U4065(__A04_NET_309, __A04_NET_316, __A04_NET_311, __A04_2__BRXP3, T03_n, IC15_n, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC4002 U4066(RSC_n, __A04_NET_315, __A04_NET_323, __A04_NET_308, __A04_2__BRXP3,  , GND,  , __A04_NET_315, __A04_NET_303, __A04_NET_323, __A04_2__BRXP3, __A04_NET_302, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5001(IC10, IC3, TC0, TCF0, IC4, __A05_NET_215, GND, __A05_NET_216, IC2, IC3, RSM3, __A05_NET_217, IC2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5002(__A05_NET_218, STD2, IC2, __A05_NET_203, T01_n, __A05_NET_217, GND, T01_n, __A05_NET_218, __A05_NET_187, IC10_n, T01_n, __A05_NET_186, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5003(__A05_NET_188, T01_n, __A05_NET_215, __A05_NET_185, T02_n, __A05_NET_216, GND, T08_n, CCS0_n, __A05_NET_257, T02_n, MP3_n, n2XP7, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U5004(T02_n, STD2, __A05_1__10XP6, __A05_1__10XP7, __A05_NET_186, __A05_NET_213, GND, __A05_NET_212, __A05_NET_187, n3XP6, __A05_NET_191, DVST, DIV_n, VCC, SIM_RST, SIM_CLK);
    assign MONEX_n = MONEX_n_U5005_2;
    assign RZ_n = RZ_n_U5005_4;
    assign RB_n = RB_n_U5005_6;
    assign RA_n = RA_n_U5005_8;
    assign WA_n = WA_n_U5005_10;
    assign RL_n = RL_n_U5005_12;
    U74LVC07 U5005(__A05_NET_213, MONEX_n_U5005_2, __A05_NET_212, RZ_n_U5005_4, __A05_NET_207, RB_n_U5005_6, GND, RA_n_U5005_8, __A05_NET_214, WA_n_U5005_10, __A05_NET_221, RL_n_U5005_12, __A05_NET_220, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5006(__A05_NET_185, __A05_1__8XP15, __A05_NET_195, __A05_NET_190, __A05_1__8XP12, __A05_NET_220, GND, __A05_1__PARTC, INKL_n, SHIFT, MONpCH, __A05_1__NISQ_n, n2XP7, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5007(__A05_1__3XP5, T03_n, IC2_n, __A05_NET_177, T01_n, IC15_n, GND, __A05_NET_177, __A05_NET_184, __A05_NET_214, T03_n, TC0_n, n3XP6, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5008(__A05_NET_184, T04_n, IC2_n, __A05_NET_193, T02_n, IC15_n, GND, __A05_NET_193, __A05_NET_178, TPZG_n, T04_n, DAS0_n, __A05_NET_195, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U5009(__A05_NET_221, __A05_NET_195, __A05_NET_194, __A05_NET_194, T04_n, MASK0_n, GND, MP3_n, T10_n, __A05_NET_190, T05_n, IC2_n, __A05_NET_191, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5010(__A05_NET_178, T05_n, __A05_NET_180, __A05_NET_219, __A05_NET_177, __A05_NET_178, GND, T05_n, DAS0_n, n5XP12, T06_n, RSM3_n, __A05_NET_209, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5011(__A05_1__PARTC, PRINC, __A05_NET_178, __A05_NET_177, n7XP9, __A05_NET_179, GND, __A05_NET_182, n9XP5, __A05_NET_177, __A05_NET_209, __A05_NET_180, CCS0, VCC, SIM_RST, SIM_CLK);
    assign TMZ_n = TMZ_n_U5012_2;
    assign WG_n = WG_n_U5012_4;
    assign RG_n = RG_n_U5012_6;
    assign RC_n = RC_n_U5012_8;
    assign A2X_n = A2X_n_U5012_10;
    assign WY_n = WY_n_U5012_12;
    U74LVC07 U5012(__A05_NET_219, TMZ_n_U5012_2, __A05_NET_182, WG_n_U5012_4, __A05_NET_181, RG_n_U5012_6, GND, RC_n_U5012_8, __A05_NET_205, A2X_n_U5012_10, __A05_NET_199, WY_n_U5012_12, __A05_NET_196, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5013(__A05_NET_197, T06_n, DAS0_n, __A05_NET_208, T06_n, MSU0_n, GND, __A05_NET_194, __A05_NET_208, __A05_NET_205, T07_n, DAS0_n, __A05_NET_206, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b1) U5014(__A05_NET_178, __A05_NET_198, __A05_NET_198, __A05_NET_197, __A05_NET_208, __A05_NET_199, GND, __A05_NET_196, __A05_NET_198, __A05_NET_208, __A05_NET_197, __A05_NET_181, __A05_NET_197, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U5015(__A05_NET_207, __A05_NET_188, __A05_1__3XP5, __A05_NET_206, __A05_NET_209,  , GND,  , IC3, RSM3, MP3, IC16, TSUDO_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5016(n7XP9, T07_n, MSU0_n, __A05_NET_198, T07_n, IC2_n, GND, T07_n, CCS0_n, __A05_NET_246, __A05_NET_243, __A05_NET_244, __A05_NET_239, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U5017(__A05_NET_208, __A05_NET_203, __A05_1__8XP3, __A05_NET_246, n4XP5, __A05_NET_202, GND, __A05_NET_247, n4XP5, __A05_NET_246, __A05_NET_203, __A05_NET_200, __A05_1__10XP6, VCC, SIM_RST, SIM_CLK);
    assign CI_n = CI_n_U5018_2;
    assign RZ_n = RZ_n_U5018_4;
    assign WY12_n = WY12_n_U5018_6;
    assign WZ_n = WZ_n_U5018_8;
    assign RB_n = RB_n_U5018_10;
    assign WB_n = WB_n_U5018_12;
    U74LVC07 U5018(__A05_NET_200, CI_n_U5018_2, __A05_NET_202, RZ_n_U5018_4, __A05_NET_247, WY12_n_U5018_6, GND, WZ_n_U5018_8, __A05_NET_242, RB_n_U5018_10, __A05_NET_239, WB_n_U5018_12, __A05_NET_245, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U5019(CCS0_n, T07_n, BR1_n, CCS0_n, T07_n, PTWOX, GND, __A05_NET_242, __A05_1__3XP5, __A05_NET_249, __A05_NET_257, n7XP4, BR2_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5020(INKL_n, FETCH0, __A05_NET_257, __A05_NET_255, n9XP5, __A05_NET_254, GND, __A05_NET_256, IC2, IC4, DXCH0, __A05_NET_243, T08_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U5021(RAD, TSUDO_n, T08_n, __A05_NET_245, RAD, __A05_NET_250, GND, T08_n, __A05_NET_253, __A05_1__8XP15, T08_n, __A05_NET_252, __A05_1__8XP3, VCC, SIM_RST, SIM_CLK);
    U74HC04 U5022(IC16, __A05_NET_253, __A05_NET_350, RQ_n, MP3, __A05_NET_263, GND, SCAD_n, SCAD, NDR100_n, __A05_NET_260, __A05_NET_321, __A05_NET_274, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5023(__A05_NET_252, MP0, IC1, __A05_NET_255, T08_n, __A05_NET_256, GND, T08_n, __A05_NET_248, __A05_NET_250, T08_n, GOJ1_n, RSTRT, VCC, SIM_RST, SIM_CLK);
    assign RU_n = RU_n_U5024_2;
    assign RA_n = RA_n_U5024_4;
    assign ST2_n = ST2_n_U5024_6;
    assign WY_n = WY_n_U5024_8;
    assign RC_n = RC_n_U5024_10;
    assign WA_n = WA_n_U5024_12;
    U74LVC07 U5024(__A05_NET_254, RU_n_U5024_2, __A05_NET_229, RA_n_U5024_4, __A05_NET_230, ST2_n_U5024_6, GND, WY_n_U5024_8, __A05_NET_222, RC_n_U5024_10, __A05_NET_236, WA_n_U5024_12, __A05_NET_233, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5025(DXCH0, GOJ1, CCS0_n, BR2, T10_n, __A05_1__10XP6, GND, __A05_NET_225, IC1, IC10, RUPT0, __A05_NET_248, DAS0, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5026(__A05_1__8XP12, T08_n, DAS0_n, __A05_NET_249, T08_n, TCSAJ3_n, GND, T09_n, __A05_NET_251, __A05_NET_244, IC2, __A05_1__DV1B1B, __A05_NET_251, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5027(n9XP5, T09_n, DAS0_n, __A05_NET_223, T09_n, MASK0_n, GND, __A05_NET_223, __A05_NET_224, __A05_NET_229, T10_n, CCS0_n, __A05_NET_231, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5028(__A05_NET_230, __A05_NET_249, __A05_NET_231, n10XP1, __A05_NET_225, T10_n, GND, T10_n, __A05_NET_228, __A05_NET_224, DAS0, __A05_NET_226, __A05_NET_228, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U5029(__A05_NET_231, __A05_NET_223, T10_n, DAS0_n, BR1B2_n, n10XP8, GND, __A05_NET_233, __A05_NET_244, __A05_NET_234, n5XP11, __A05_NET_222, __A05_NET_224, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5030(__A05_NET_226, MSU0_n, BR1_n, __A05_1__10XP7, T10_n, __A05_NET_227, GND, __A05_NET_226, __A05_NET_235, __A05_NET_227, BR12B_n, DAS0_n, __A05_NET_235, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5031(n11XP2, T11_n, MSU0_n, __A05_NET_238, T11_n, MASK0_n, GND, __A05_NET_223, __A05_NET_238, __A05_NET_236, T11_n, __A05_NET_237, __A05_NET_234, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5032(__A05_NET_237, MSU0, IC14,  ,  ,  , GND, GOJAM, GNHNC, __A05_NET_232, __A05_NET_232, T01, GNHNC, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U5034( ,  , IC12, DAS0, DAS1, __A05_NET_297, GND, __A05_NET_304, RL10BB, __A05_NET_302, RSCT,  ,  , VCC, SIM_RST, SIM_CLK);
    assign __A05_NET_299 = __A05_NET_299_U5035_8;
    assign __A05_NET_299 = __A05_NET_299_U5035_10;
    assign WS_n = WS_n_U5035_12;
    U74LVC07 U5035( ,  ,  ,  ,  ,  , GND, __A05_NET_299_U5035_8, __A05_NET_297, __A05_NET_299_U5035_10, __A05_NET_298, WS_n_U5035_12, __A05_NET_304, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5036( ,  ,  ,  ,  ,  , GND, T01_n, __A05_NET_299, RL10BB, T01_n, FETCH0_n, R6, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U5037(__A05_NET_298, IC9, DXCH0, PRINC, INOUT,  , GND,  , YB0_n, YT0_n, S12, S11, __A05_NET_260, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5038(__A05_NET_302, T01_n, CHINC_n, __A05_NET_351, T03_n, __A05_NET_303, GND, IC5, MP0, __A05_NET_293, T03_n, IC8_n, __A05_NET_296, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U5039(T01_n, MONpCH, TS0, DAS0, MASK0, __A05_NET_294, GND, __A05_NET_291, __A05_NET_351, __A05_NET_296, __A05_NET_350, RSCT, INKL_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U5040(__A05_NET_314, __A05_NET_349,  ,  ,  ,  , GND,  ,  ,  ,  , __A05_NET_292, __A05_2__6XP2, VCC, SIM_RST, SIM_CLK);
    assign WB_n = WB_n_U5041_2;
    assign WB_n = WB_n_U5041_4;
    assign __A05_NET_303 = __A05_NET_303_U5041_6;
    assign __A05_NET_303 = __A05_NET_303_U5041_8;
    assign RL_n = RL_n_U5041_10;
    assign RA_n = RA_n_U5041_12;
    U74LVC07 U5041(__A05_NET_291, WB_n_U5041_2, __A05_NET_292, WB_n_U5041_4, __A05_NET_294, __A05_NET_303_U5041_6, GND, __A05_NET_303_U5041_8, __A05_NET_293, RL_n_U5041_10, __A05_NET_295, RA_n_U5041_12, __A05_NET_315, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5042(n2XP8, T02_n, FETCH0_n, __A05_NET_350, T03_n, QXCH0_n, GND, T04_n, DV1_n, __A05_NET_316, T04_n, __A05_NET_320, __A05_NET_314, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5043(__A05_NET_296, __A05_NET_316, DV1, INOUT, IC2, __A05_NET_320, GND, __A05_NET_317, __A05_NET_349, __A05_NET_309, __A05_2__5XP9, __A05_NET_295, __A05_2__11XP6, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5044(__A05_NET_315, __A05_NET_351, __A05_2__6XP2, TRSM, T05_n, NDX0_n, GND, IC12_n, T05_n, __A05_NET_349, DAS1_n, T05_n, __A05_NET_309, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U5045(__A05_2__5XP13, n5XP15, DAS1, PRINC, __A05_1__PARTC, __A05_NET_310, GND, __A05_NET_306, __A05_NET_308, n2XP8, __A05_2__10XP10, __A05_NET_319, __A05_NET_347, VCC, SIM_RST, SIM_CLK);
    assign RG_n = RG_n_U5046_2;
    assign RG_n = RG_n_U5046_4;
    assign WY_n = WY_n_U5046_6;
    assign A2X_n = A2X_n_U5046_8;
    assign CI_n = CI_n_U5046_10;
    assign WY12_n = WY12_n_U5046_12;
    U74LVC07 U5046(__A05_NET_317, RG_n_U5046_2, __A05_NET_319, RG_n_U5046_4, __A05_NET_306, WY_n_U5046_6, GND, A2X_n_U5046_8, __A05_NET_307, CI_n_U5046_10, __A05_NET_311, WY12_n_U5046_12, __A05_NET_265, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U5047(__A05_NET_308, __A05_NET_310, T05_n, __A05_NET_307, __A05_NET_309, __A05_2__10XP10, GND, SHIFT_n, T05_n, __A05_2__5XP9, SHANC_n, T05_n, __A05_NET_313, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5048(__A05_NET_313, __A05_NET_346, YT0_n, YB0_n, XT0_n, __A05_NET_262, GND, __A05_NET_282, RAND0, WAND0, __A05_NET_274, __A05_NET_311, __A05_NET_264, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5049(__A05_2__5XP13, IC8_n, T05_n, n5XP15, QXCH0_n, T05_n, GND, CHINC_n, T05_n, n5XP21, IC5_n, T05_n, __A05_NET_347, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U5050(__A05_NET_346, IC16_n, T05_n, __A05_NET_264, __A05_NET_263, T05_n, GND, __A05_NET_346, __A05_NET_264, __A05_NET_265, S11, S12, __A05_NET_261, VCC, SIM_RST, SIM_CLK);
    assign RB_n = RB_n_U5051_2;
    assign RZ_n = RZ_n_U5051_4;
    assign SCAD = SCAD_U5051_6;
    assign SCAD = SCAD_U5051_8;
    assign RC_n = RC_n_U5051_10;
    assign __A05_NET_287 = __A05_NET_287_U5051_12;
    U74LVC07 U5051(__A05_NET_268, RB_n_U5051_2, __A05_NET_266, RZ_n_U5051_4, __A05_NET_261, SCAD_U5051_6, GND, SCAD_U5051_8, __A05_NET_262, RC_n_U5051_10, __A05_NET_279, __A05_NET_287_U5051_12, __A05_NET_288, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5052(__A05_NET_268, __A05_2__5XP19, __A05_NET_346, __A05_NET_266, __A05_2__6XP7, __A05_NET_264, GND, XT2_n, NDR100_n, OCTAD2, NDR100_n, XT3_n, OCTAD3, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5053(OCTAD4, NDR100_n, XT4_n, OCTAD5, NDR100_n, XT5_n, GND, NDR100_n, XT6_n, OCTAD6, BR1_n, DV1_n, __A05_NET_274, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5054(__A05_NET_283, __A05_NET_282, T05_n, __A05_2__5XP19, T05_n, __A05_NET_281, GND, DV1_n, BR1, __A05_1__DV1B1B, TS0_n, BRDIF_n, __A05_NET_290, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b0, 1'b1) U5055(__A05_NET_279, __A05_NET_283, __A05_NET_284, __A05_NET_339, __A05_NET_285,  , GND,  , __A05_2__5XP13, __A05_NET_337, __A05_NET_326, __A05_NET_332, __A05_NET_327, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5056(ROR0, __A05_1__DV1B1B, IC2, IC5, READ0, __A05_NET_288, GND, __A05_NET_277, IC2, IC3, TS0, __A05_NET_281, WOR0, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U5057(__A05_NET_289, __A05_NET_290, DV4, __A05_NET_272, __A05_NET_287, T05_n, GND, __A05_NET_321, T05_n, __A05_NET_273, __A05_NET_272, __A05_NET_284, __A05_NET_271, VCC, SIM_RST, SIM_CLK);
    assign __A05_NET_287 = __A05_NET_287_U5058_2;
    assign Z16_n = Z16_n_U5058_4;
    assign WA_n = WA_n_U5058_6;
    assign __A05_NET_278 = __A05_NET_278_U5058_8;
    assign __A05_NET_278 = __A05_NET_278_U5058_10;
    assign WZ_n = WZ_n_U5058_12;
    U74LVC07 U5058(__A05_NET_289, __A05_NET_287_U5058_2, __A05_NET_270, Z16_n_U5058_4, __A05_NET_271, WA_n_U5058_6, GND, __A05_NET_278_U5058_8, __A05_NET_277, __A05_NET_278_U5058_10, __A05_NET_275, WZ_n_U5058_12, __A05_NET_276, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0) U5059(__A05_NET_273, __A05_NET_270, __A05_NET_330, __A05_NET_276, __A05_NET_284, __A05_NET_322, GND, __A05_NET_338, __A05_NET_339, NISQ, __A05_1__NISQ_n, __A05_1__MNISQ, __A05_1__NISQ_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U5060(__A05_NET_275, IC16, MP3, __A05_NET_330, T06_n, __A05_NET_278, GND, T06_n, DAS1_n, n6XP8, n6XP8, __A05_2__6XP7, __A05_NET_345, VCC, SIM_RST, SIM_CLK);
    assign TOV_n = TOV_n_U5061_2;
    assign RU_n = RU_n_U5061_4;
    assign RU_n = RU_n_U5061_6;
    assign WB_n = WB_n_U5061_8;
    assign RG_n = RG_n_U5061_10;
    assign TSGN_n = TSGN_n_U5061_12;
    U74LVC07 U5061(__A05_NET_345, TOV_n_U5061_2, __A05_NET_343, RU_n_U5061_4, __A05_NET_344, RU_n_U5061_6, GND, WB_n_U5061_8, __A05_NET_341, RG_n_U5061_10, __A05_NET_342, TSGN_n_U5061_12, __A05_NET_323, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5062(__A05_2__6XP7, DV4_n, T06_n, __A05_NET_329, T07_n, __A05_NET_331, GND, T07_n, STFET1_n, __A05_NET_328, T08_n, DV4_n, RSTSTG, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5063(__A05_NET_330, n6XP8, __A05_NET_336, __A05_NET_326, __A05_NET_337, __A05_NET_344, GND, __A05_2__6XP2, T06_n, RXOR0, INOUT_n, __A05_NET_343, n5XP11, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U5064(IC13, IC14, __A05_NET_329, __A05_NET_326, __A05_NET_336, __A05_NET_341, GND, __A05_NET_342, __A05_NET_329, __A05_NET_328, __A05_NET_285, __A05_NET_331, DV1, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5065(T08_n, MONWBK, IC2, IC14, DV1, __A05_NET_335, GND, __A05_NET_333, DV4B1B, IC4, __A05_NET_334, U2BBK, STFET1_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U5066(__A05_NET_323, RSTSTG, __A05_2__5XP9, __A05_NET_284, T09_n, __A05_NET_321, GND, T09_n, DV4_n, __A05_NET_326, T09_n, DAS1_n, __A05_NET_339, VCC, SIM_RST, SIM_CLK);
    assign Z15_n = Z15_n_U5067_2;
    assign WL_n = WL_n_U5067_4;
    assign TMZ_n = TMZ_n_U5067_6;
    assign WYD_n = WYD_n_U5067_8;
    assign TSGN_n = TSGN_n_U5067_10;
    U74LVC07 U5067(__A05_NET_322, Z15_n_U5067_2, __A05_NET_327, WL_n_U5067_4, __A05_NET_338, TMZ_n_U5067_6, GND, WYD_n_U5067_8, __A05_NET_340, TSGN_n_U5067_10, __A05_NET_179,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U5068(__A05_NET_336, T10_n, __A05_NET_335,  ,  ,  , GND, T10_n, IC11_n, __A05_2__10XP10, T10_n, __A05_NET_333, __A05_NET_332, VCC, SIM_RST, SIM_CLK);
    U74HC27 U5069(DAS1_n, ADS0, T12_n, T12USE_n, DV1_n, __A05_NET_337, GND,  ,  ,  ,  , __A05_NET_334, BR2, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U5070(DV4B1B, DV4_n, BR1, __A05_2__11XP6, T11_n, DV1_n, GND, __A05_2__5XP9, __A05_2__11XP6, __A05_NET_340, T11_n, RXOR0_n, __A05_NET_285, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6001(T04, T07, __A06_NET_288, __A06_NET_289, __A06_NET_290, __A06_NET_287, GND, __A06_NET_305, T01, T03, T05, __A06_NET_302, T10, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6002(__A06_NET_288, __A06_NET_302, DV376_n, __A06_NET_289, T01_n, DV1376_n, GND, T04_n, DV4_n, __A06_NET_290, MP1_n, __A06_NET_291, __A06_NET_292, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U6003(T07, T09, __A06_1__L15A_n, __A06_1__L02A_n, L01_n, __A06_NET_304, GND, __A06_NET_345, T05, T08, T11, __A06_NET_306, T11, VCC, SIM_RST, SIM_CLK);
    assign __A06_NET_291 = __A06_NET_291_U6004_2;
    assign __A06_NET_291 = __A06_NET_291_U6004_4;
    assign A2X_n = A2X_n_U6004_6;
    assign RB_n = RB_n_U6004_8;
    assign WYD_n = WYD_n_U6004_10;
    assign WY_n = WY_n_U6004_12;
    U74LVC07 U6004(__A06_NET_305, __A06_NET_291_U6004_2, __A06_NET_306, __A06_NET_291_U6004_4, __A06_NET_303, A2X_n_U6004_6, GND, RB_n_U6004_8, __A06_NET_317, WYD_n_U6004_10, __A06_NET_318, WY_n_U6004_12, __A06_NET_309, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b0) U6005(__A06_NET_316, __A06_NET_292, n2XP7, L2GD_n, __A06_1__ZIP, __A06_1__DVXP1, GND, __A06_1__DVXP1, __A06_NET_310, __A06_NET_318, __A06_NET_307, __A06_NET_308, __A06_NET_311, VCC, SIM_RST, SIM_CLK);
    U74HC04 U6006(L01_n, __A06_NET_294, __A06_1__L02A_n, __A06_NET_344, __A06_1__L15A_n, __A06_NET_293, GND, __A06_1__DVXP1, __A06_NET_287, __A06_1__ZIP, __A06_NET_316, __A06_NET_342, __A06_NET_343, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U6007(n7XP19, __A06_1__ZIP, __A06_1__DVXP1, __A06_NET_313, RBSQ, __A06_NET_317, GND, __A06_NET_320, __A06_NET_294, __A06_NET_344, __A06_NET_293, __A06_NET_303, __A06_1__DVXP1, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6008(__A06_NET_293, __A06_NET_294, __A06_NET_316, __A06_NET_308, __A06_NET_307, __A06_NET_319, GND, __A06_NET_343, __A06_NET_307, __A06_NET_308, __A06_1__L02A_n, __A06_NET_308, __A06_1__L02A_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6009(__A06_NET_310, __A06_NET_316, __A06_NET_311, __A06_NET_315, __A06_NET_316, __A06_NET_342, GND, __A06_NET_345, DV376_n, __A06_NET_314, DV1376_n, T02_n, __A06_NET_276, VCC, SIM_RST, SIM_CLK);
    U74HC04 U6010(__A06_NET_315, MCRO_n, __A06_NET_281, __A06_NET_278, __A06_NET_285, __A06_NET_286, GND, __A06_1__ZAP, ZAP_n, __A06_NET_347, __A06_NET_345, MONEX, MONEX_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6011(__A06_NET_316, __A06_NET_342, __A06_NET_343, __A06_NET_320, __A06_NET_316, __A06_NET_313, GND, __A06_NET_307, __A06_NET_344, __A06_1__L15A_n, L01_n, __A06_1__ZIPCI, __A06_NET_304, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b0) U6012(__A06_NET_281, __A06_NET_314, __A06_NET_276, __A06_NET_285, __A06_NET_280, DIVSTG, GND, T08, T10, __A06_NET_282, MP1_n, __A06_NET_284, __A06_NET_270, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U6013(T06, T09, DV376_n, __A06_NET_279, T12USE_n, __A06_NET_280, GND, __A06_NET_283, T02, T04, T06, __A06_NET_279, T12, VCC, SIM_RST, SIM_CLK);
    assign __A06_NET_284 = __A06_NET_284_U6014_2;
    assign __A06_NET_284 = __A06_NET_284_U6014_4;
    assign WL_n = WL_n_U6014_6;
    assign RG_n = RG_n_U6014_8;
    assign WB_n = WB_n_U6014_10;
    assign RU_n = RU_n_U6014_12;
    U74LVC07 U6014(__A06_NET_283, __A06_NET_284_U6014_2, __A06_NET_282, __A06_NET_284_U6014_4, __A06_NET_277, WL_n_U6014_6, GND, RG_n_U6014_8, __A06_NET_274, WB_n_U6014_10, __A06_NET_295, RU_n_U6014_12, __A06_NET_296, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U6015(__A06_NET_272, T01, T03, __A06_NET_271, __A06_NET_272, MP3_n, GND, __A06_NET_270, __A06_NET_271, ZAP_n, n5XP28, __A06_NET_278, TSGU_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b1) U6016(__A06_NET_277, __A06_NET_278, n5XP12, __A06_NET_301, RRPA, n5XP4, GND, n5XP15, n3XP6, WQ_n, n9XP5, n6XP8, __A06_NET_350, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b0, 1'b1) U6017(__A06_NET_274, n5XP4, RADRG, __A06_NET_278, n5XP28,  , GND,  , n5XP28, n1XP10, __A06_NET_286, n2XP3, __A06_NET_295, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U6018(__A06_NET_296, __A06_NET_286, __A06_1__ZAP, n5XP12, n6XP5,  , GND,  , PRINC, PINC, MINC, DINC, __A06_NET_235, VCC, SIM_RST, SIM_CLK);
    assign WZ_n = WZ_n_U6019_2;
    assign TOV_n = TOV_n_U6019_4;
    assign WSC_n = WSC_n_U6019_6;
    assign WG_n = WG_n_U6019_8;
    assign __A06_NET_268 = __A06_NET_268_U6019_10;
    assign __A06_NET_268 = __A06_NET_268_U6019_12;
    U74LVC07 U6019(__A06_NET_301, WZ_n_U6019_2, __A06_NET_349, TOV_n_U6019_4, __A06_NET_350, WSC_n_U6019_6, GND, WG_n_U6019_8, __A06_NET_346, __A06_NET_268_U6019_10, __A06_NET_269, __A06_NET_268_U6019_12, __A06_NET_219, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U6020(n6XP5, n3XP2, BR1_n, PHS4_n, TSGU_n, RB1F, GND, CLXC, TSGU_n, BR1, PHS4_n, __A06_NET_349, n9XP5, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b1) U6021(__A06_NET_346, n6XP8, n6XP8, PIFL_n, __A06_1__DVXP1, __A06_NET_348, GND, PTWOX, MONEX, __A06_NET_332, MONEX, B15X, __A06_NET_333, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U6022(PIFL_n, __A06_NET_347, STBE, n1XP10, STBF, __A06_NET_331, GND, __A06_NET_269, __A06_NET_266, __A06_NET_265, INCR0, __A06_NET_348, T02, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0) U6023(__A06_NET_332, TWOX, __A06_NET_333, BXVX, __A06_NET_324, __A06_NET_321, GND, __A06_NET_322, __A06_NET_321, __A06_NET_330, __A06_NET_322, __A06_NET_329, __A06_NET_330, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U6024(CGMC, __A06_NET_331, __A06_NET_325, __A06_NET_323, CGMC, __A06_NET_324, GND, __A06_NET_323, __A06_NET_331, __A06_NET_324, BR1, AUG0_n, __A06_NET_266, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0) U6025(__A06_NET_329, __A06_NET_328, __A06_NET_328, __A06_NET_326, __A06_NET_326, __A06_NET_327, GND, __A06_NET_325, __A06_NET_327, __A06_NET_212, __A06_NET_223, __A06_NET_239, __A06_2__7XP10, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6026(__A06_NET_265, DIM0_n, BR12B_n, __A06_NET_219, PINC, __A06_NET_267, GND, BR12B_n, DINC_n, __A06_NET_267, T06_n, __A06_NET_268, __A06_2__6XP10, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6027(__A06_NET_218, MINC, MCDU, __A06_NET_225, AUG0_n, BR1_n, GND, DIM0_n, BR1B2B_n, __A06_NET_221, BR1B2B_n, DINC_n, __A06_NET_222, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6028(__A06_NET_225, __A06_NET_221, BR1B2B_n, CDUSTB_n, DINC_n, __A06_2__POUT, GND, __A06_2__MOUT, BR12B_n, CDUSTB_n, DINC_n, __A06_NET_217, __A06_NET_222, VCC, SIM_RST, SIM_CLK);
    assign __A06_NET_224 = __A06_NET_224_U6029_2;
    assign __A06_NET_224 = __A06_NET_224_U6029_4;
    assign MONEX_n = MONEX_n_U6029_6;
    assign WA_n = WA_n_U6029_8;
    assign RB1_n = RB1_n_U6029_10;
    assign R1C_n = R1C_n_U6029_12;
    U74LVC07 U6029(__A06_NET_218, __A06_NET_224_U6029_2, __A06_NET_217, __A06_NET_224_U6029_4, __A06_NET_212, MONEX_n_U6029_6, GND, WA_n_U6029_8, __A06_NET_214, RB1_n_U6029_10, __A06_NET_239, R1C_n_U6029_12, __A06_NET_227, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6030(__A06_NET_223, T06_n, __A06_NET_224, __A06_NET_213, PCDU, MCDU, GND, T06_n, __A06_NET_213, __A06_2__6XP12, __A06_NET_216, T07_n, __A06_NET_215, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b1) U6031(BR2_n, DINC_n, DAS0, DAS1, MSU0, __A06_NET_216, GND, __A06_NET_214, __A06_NET_215, __A06_2__7XP7, __A06_NET_231, __A06_2__ZOUT, CDUSTB_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6032(__A06_NET_237, DV4_n, BR1B2B, __A06_2__7XP7, T07_n, __A06_NET_238, GND, WAND0, INOTLD, __A06_NET_241, T07_n, __A06_NET_241, n7XP14, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6033(__A06_NET_237, WAND0, DAS1_n, T07_n, BR1B2_n, __A06_2__7XP10, GND, __A06_2__7XP11, DAS1_n, T07_n, BR12B_n, __A06_NET_238, RAND0, VCC, SIM_RST, SIM_CLK);
    U74HC04 U6034(__A06_2__7XP11, __A06_NET_227, __A06_NET_199, PONEX, ST2_n, ST2, GND, ST1, __A06_NET_245, __A06_NET_250, PSEUDO, __A06_NET_249, __A06_2__RDBANK, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6035(__A06_2__7XP15, __A06_NET_226, T07_n, __A06_NET_230, __A06_NET_235, T07_n, GND, PRINC, INKL, __A06_NET_192, IC9, DXCH0, __A06_NET_193, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6036(PCDU, MCDU, n7XP9, n11XP2, __A06_2__7XP15, RUS_n, GND, __A06_NET_229, __A06_NET_230, __A06_NET_228, __A06_NET_231, __A06_NET_226, SHIFT, VCC, SIM_RST, SIM_CLK);
    assign RU_n = RU_n_U6037_2;
    assign WSC_n = WSC_n_U6037_4;
    assign WG_n = WG_n_U6037_6;
    assign RB_n = RB_n_U6037_8;
    assign n8PP4 = n8PP4_U6037_10;
    assign n8PP4 = n8PP4_U6037_12;
    U74LVC07 U6037(__A06_NET_229, RU_n_U6037_2, __A06_NET_188, WSC_n_U6037_4, __A06_NET_195, WG_n_U6037_6, GND, RB_n_U6037_8, __A06_NET_183, n8PP4_U6037_10, __A06_NET_184, n8PP4_U6037_12, __A06_NET_181, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U6038(__A06_NET_192, T07_n, T04_n, MON_n, FETCH1, __A06_NET_190, GND, __A06_NET_188, __A06_NET_189, __A06_NET_190, __A06_NET_191, __A06_NET_189, MONpCH, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6039(__A06_NET_195, __A06_NET_189, __A06_NET_191, __A06_NET_191, T07_n, __A06_NET_193, GND, __A06_2__10XP9, __A06_NET_191, __A06_NET_183, T08_n, n8PP4, __A06_2__8XP4, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6040(RUPT1, DAS1, IC17, MASK0, IC11, __A06_NET_181, GND, __A06_NET_182, IC6, IC7, IC9, __A06_NET_184, MSU0, VCC, SIM_RST, SIM_CLK);
    assign n8PP4 = n8PP4_U6041_2;
    assign __A06_NET_209 = __A06_NET_209_U6041_4;
    assign __A06_NET_209 = __A06_NET_209_U6041_6;
    assign WS_n = WS_n_U6041_8;
    assign __A06_NET_210 = __A06_NET_210_U6041_10;
    assign __A06_NET_210 = __A06_NET_210_U6041_12;
    U74LVC07 U6041(__A06_NET_182, n8PP4_U6041_2, __A06_NET_185, __A06_NET_209_U6041_4, __A06_NET_186, __A06_NET_209_U6041_6, GND, WS_n_U6041_8, __A06_NET_204, __A06_NET_210_U6041_10, __A06_NET_206, __A06_NET_210_U6041_12, __A06_NET_205, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U6042(T08_n, RUPT0, __A06_NET_209, R6, R15, __A06_NET_204, GND, __A06_NET_205, ADS0, IC11, __A06_NET_207, __A06_NET_185, DAS0, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6043(__A06_NET_186, MP1, DV1376, __A06_NET_208, MP3_n, BR1_n, GND, __A06_NET_208, CCS0, __A06_NET_206, T11_n, __A06_NET_210, __A06_NET_231, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6044(__A06_NET_207, DAS1_n, BR2_n, __A06_NET_198, __A06_1__ZIPCI, __A06_2__6XP12, GND, CCS0_n, BR1B2B_n, __A06_NET_201, T10_n, NDXX1_n, EXT, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U6045(T03_n, DAS1_n, __A06_NET_243, __A06_NET_228, n2XP5, __A06_NET_262, GND, __A06_NET_264, IC7, DCS0, SU0, __A06_NET_228, ADS0, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U6046(__A06_NET_199, n8XP6, n7XP4, n10XP8, __A06_2__6XP10,  , GND,  , IC6, DCA0, AD0, __A06_NET_201, __A06_NET_200, VCC, SIM_RST, SIM_CLK);
    assign CI_n = CI_n_U6047_2;
    assign WA_n = WA_n_U6047_4;
    assign RC_n = RC_n_U6047_6;
    assign __A06_NET_248 = __A06_NET_248_U6047_8;
    assign __A06_NET_248 = __A06_NET_248_U6047_10;
    assign ST2_n = ST2_n_U6047_12;
    U74LVC07 U6047(__A06_NET_198, CI_n_U6047_2, __A06_NET_262, WA_n_U6047_4, __A06_NET_263, RC_n_U6047_6, GND, __A06_NET_248_U6047_8, __A06_NET_264, __A06_NET_248_U6047_10, __A06_NET_259, ST2_n_U6047_12, __A06_NET_258, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6048(__A06_2__10XP9, T10_n, __A06_NET_200, __A06_NET_244, IC6, IC7, GND, T10_n, __A06_NET_244, __A06_NET_243, T10_n, __A06_NET_248, __A06_NET_247, VCC, SIM_RST, SIM_CLK);
    U74HC02 U6049(__A06_NET_263, __A06_NET_247, __A06_2__7XP7, __A06_NET_259, __A06_NET_246, DV4B1B, GND, CCS0_n, BR12B_n, __A06_NET_246, T10_n, MP1_n, __A06_2__10XP15, VCC, SIM_RST, SIM_CLK);
    U74HC27 U6050(__A06_2__8XP4, __A06_2__10XP15, __A06_2__8XP4, RADRZ, n9XP1, __A06_NET_256, GND, NEAC, __A06_NET_255, TL15, GOJAM, __A06_NET_258, RADRZ, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U6051(__A06_NET_245, n2XP8, n10XP1, MP0T10, __A06_2__10XP15,  , GND,  , __A06_1__DVXP1, GOJAM, NISQ, __A06_1__WHOMP_n, WHOMP, VCC, SIM_RST, SIM_CLK);
    assign RZ_n = RZ_n_U6052_2;
    assign RPTSET = RPTSET_U6052_4;
    assign RU_n = RU_n_U6052_6;
    assign RC_n = RC_n_U6052_8;
    U74LVC07 U6052(__A06_NET_256, RZ_n_U6052_2, __A06_NET_250, RPTSET_U6052_4, __A06_NET_249, RU_n_U6052_6, GND, RC_n_U6052_8, __A06_NET_340,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U6053(__A06_NET_255, MP0T10, NEAC, __A06_NET_257, RADRZ, PSEUDO, GND, T06_n, STFET1_n, __A06_2__RDBANK, __A06_1__ZIPCI, n3XP7, __A06_NET_340, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U6054(__A06_NET_257, GOJAM, n3XP7, n5XP21, n4XP11, RCH_n, GND,  ,  ,  ,  , PSEUDO, RADRG, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U6055(R1C_n, R1C, RB1_n, RB1, L02_n, __A06_NET_334, GND, __A06_1__L02A_n, __A06_NET_334, __A06_NET_335, L15_n, __A06_1__L15A_n, __A06_NET_335, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U6056(__A06_NET_319, __A06_NET_309, __A06_1__WHOMP_n, WHOMPA, __A06_NET_189, WOVR_n, GND, POUT_n, __A06_2__POUT, MOUT_n, __A06_2__MOUT, ZOUT_n, __A06_2__ZOUT, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U6057(__A06_1__WHOMP_n, WHOMP, CLXC,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U7001(__A07_1__WALSG, ZAP_n, WT_n, __A07_NET_166, __A07_NET_165, __A07_NET_167, GND, __A07_NET_166, WT_n, __A07_NET_169, WY_n, WT_n, __A07_NET_168, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0) U7002(__A07_1__WALSG, WALSG_n, WY12_n, __A07_NET_165, WY_n, __A07_NET_167, GND, WYLOG_n, __A07_NET_169, WYHIG_n, __A07_NET_168, __A07_1__MWYG, __A07_NET_160, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U7003(__A07_NET_160, __A07_NET_169, __A07_NET_158, __A07_NET_158, WYD_n, WT_n, GND, __A07_NET_160, CT_n, CUG, L15_n, PIFL_n, __A07_NET_164, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1) U7004(__A07_NET_158, WYDG_n, __A07_NET_162, WYDLOG_n, __A07_NET_163, WBG_n, GND, __A07_1__MWBG, WBG_n, __A07_1__MWG, __A07_1__WGA_n, WG1G_n, __A07_1__WGNORM, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U7005(__A07_NET_159, WYD_n, WT_n, __A07_NET_163, WB_n, WT_n, GND, WBG_n, CT_n, CBG, __A07_1__WGNORM, __A07_NET_175, WG2G_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U7006(SHIFT, NEAC, __A07_1__WGA_n, WT_n, GINH, __A07_1__WGNORM, GND, __A07_NET_175, __A07_1__WGA_n, WT_n, SR_n, __A07_NET_161, __A07_NET_164, VCC, SIM_RST, SIM_CLK);
    assign __A07_NET_162 = __A07_NET_162_U7007_2;
    assign __A07_NET_162 = __A07_NET_162_U7007_4;
    U74LVC07 U7007(__A07_NET_159, __A07_NET_162_U7007_2, __A07_NET_161, __A07_NET_162_U7007_4,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U7008(__A07_1__WGA_n, WT_n, __A07_1__WGA_n, WT_n, CYL_n, __A07_NET_170, GND, __A07_NET_174, __A07_1__WGA_n, WT_n, EDOP_n, __A07_NET_171, CYR_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U7009(__A07_NET_171, WG5G_n, __A07_NET_170, WG3G_n, __A07_NET_174, WEDOPG_n, GND, __A07_1__MWZG, WZG_n, __A07_1__MWLG, WLG_n, __A07_1__MWAG, WAG_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U7010(WG4G_n, __A07_NET_175, __A07_NET_171, __A07_NET_172, WT_n, WZ_n, GND, __A07_1__WSCG_n, XB5_n, __A07_NET_173, __A07_NET_172, __A07_NET_173, WZG_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7011(CZG, WZG_n, CT_n, __A07_NET_142, WL_n, WT_n, GND, __A07_1__WSCG_n, XB1_n, __A07_NET_145, __A07_NET_138, CT_n, CLG1G, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U7012(XB1_n, XT0_n, __A07_NET_142, __A07_NET_148, __A07_NET_145, WLG_n, GND, __A07_NET_139, __A07_NET_140, __A07_NET_141, __A07_1__WALSG, __A07_NET_148, WCHG_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U7013(__A07_NET_137, __A07_NET_142, __A07_NET_148, __A07_NET_145, __A07_1__WALSG,  , GND,  , __A07_NET_145, __A07_NET_148, __A07_NET_142, __A07_2__G2LSG, __A07_NET_138, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U7014(CLG2G, __A07_NET_137, CT_n, __A07_NET_140, WT_n, WA_n, GND, __A07_1__WSCG_n, XB0_n, __A07_NET_141, __A07_NET_140, __A07_NET_141, WAG_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7015(CAG, __A07_NET_139, CT_n, __A07_NET_155, WT_n, WS_n, GND, WSG_n, CT_n, CSG, WT_n, WQ_n, __A07_NET_154, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1) U7016(__A07_NET_155, WSG_n, WSG_n, __A07_1__MWSG, WQG_n, __A07_1__MWQG, GND, __A07_1__P04A, P04_n, RCG_n, __A07_NET_210, G2LSG_n, __A07_2__G2LSG, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U7017(__A07_NET_154, __A07_NET_157, XB2_n, XT0_n, WCHG_n, __A07_NET_156, GND, __A07_1__PIPSAM_n, PIPPLS_n, SB2_n, __A07_1__P04A, WQG_n, __A07_NET_156, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7018(__A07_NET_157, __A07_1__WSCG_n, XB2_n, CQG, WQG_n, CT_n, GND, RT_n, RC_n, __A07_NET_210, RT_n, RQ_n, __A07_NET_211, VCC, SIM_RST, SIM_CLK);
    U74HC27 U7019(__A07_NET_211, __A07_NET_208, XB2_n, XT0_n, __A07_2__RCHG_n, __A07_NET_209, GND, RFBG_n, __A07_NET_213, __A07_NET_215, __A07_2__RBBK, RQG_n, __A07_NET_209, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7020(__A07_NET_208, __A07_2__RSCG_n, XB2_n, __A07_NET_213, __A07_2__RSCG_n, XB4_n, GND, __A07_2__RSCG_n, XB6_n, __A07_NET_215, __A07_NET_215, __A07_2__RBBK, RBBEG_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7021(__A07_2__G2LSG, TT_n, ZAP_n, __A07_NET_212, TT_n, L2GD_n, GND, TT_n, A2X_n, __A07_NET_205, T10_n, STFET1_n, __A07_2__RBBK, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1) U7022(__A07_NET_212, L2GDG_n, __A07_NET_205, A2XG_n, __A07_NET_207, CGG, GND, __A07_2__MWEBG, WEBG_n, __A07_2__MWFBG, WFBG_n, WBBEG_n, __A07_NET_184, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7023(__A07_NET_204, L2GD_n, CT_n, __A07_NET_206, CT_n, WG_n, GND, __A07_1__WSCG_n, XB3_n, __A07_NET_185, __A07_NET_186, CT_n, CEBG, VCC, SIM_RST, SIM_CLK);
    U74HC27 U7024(__A07_NET_204, __A07_NET_206, __A07_NET_185, U2BBK, __A07_NET_184, __A07_NET_186, GND, __A07_NET_187, __A07_NET_184, U2BBK, __A07_NET_183, __A07_NET_207, CGMC, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U7025(CFBG, __A07_NET_187, CT_n, __A07_NET_183, __A07_1__WSCG_n, XB4_n, GND, __A07_NET_183, __A07_NET_184, WFBG_n, __A07_1__WSCG_n, XB6_n, __A07_NET_184, VCC, SIM_RST, SIM_CLK);
    U74HC04 U7026(WBBEG_n, __A07_2__MWBBEG, __A07_NET_191, RGG_n, RGG_n, __A07_2__MRGG, GND, __A07_2__MRAG, RAG_n, __A07_2__MRLG, RLG_n, REBG_n, __A07_NET_181, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7027(__A07_NET_191, RT_n, RG_n, __A07_NET_190, RT_n, RA_n, GND, __A07_NET_190, __A07_NET_192, RAG_n, XB0_n, __A07_2__RSCG_n, __A07_NET_192, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7028(__A07_NET_188, RT_n, RL_n, __A07_NET_189, __A07_2__RSCG_n, XB1_n, GND, RT_n, RZ_n, __A07_NET_179, __A07_NET_179, __A07_NET_177, RZG_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U7029(__A07_NET_188, __A07_NET_189, XB1_n, XT0_n, __A07_2__RCHG_n, __A07_NET_178, GND, US2SG, __A07_2__RUSG_n, SUMA15_n, SUMB15_n, RLG_n, __A07_NET_178, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7030(__A07_NET_177, XB5_n, __A07_2__RSCG_n, __A07_NET_181, __A07_2__RSCG_n, XB3_n, GND, RT_n, RU_n, __A07_NET_182, RT_n, RUS_n, __A07_NET_180, VCC, SIM_RST, SIM_CLK);
    U74HC04 U7031(__A07_NET_182, RUG_n, __A07_NET_180, __A07_2__RUSG_n, RULOG_n, __A07_2__MRULOG, GND, RBHG_n, __A07_NET_203, __A07_NET_198, RL10BB,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U7032(RULOG_n, __A07_NET_182, __A07_NET_180, __A07_NET_203, RT_n, RB_n, GND, RT_n, __A07_NET_198, __A07_NET_199, __A07_NET_203, __A07_NET_199, RBLG_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0) U7037(__A07_NET_185, WEBG_n,  ,  ,  ,  , GND, __A07_NET_202, CI_n, __A07_1__WSCG_n, __A07_NET_149, __A07_2__RSCG_n, __A07_NET_194, VCC, SIM_RST, SIM_CLK);
    U74HC27 U7038( ,  , NEAC, EAC_n, MP3A, __A07_2__CINORM, GND, __A07_NET_194, RT_n, RSC_n, SCAD_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U7039(__A07_NET_201, __A07_NET_202, __A07_2__CIFF, __A07_2__CIFF, __A07_NET_201, CUG, GND, __A07_2__CIFF, __A07_2__CINORM, CI01_n, WSC_n, SCAD_n, __A07_NET_149, VCC, SIM_RST, SIM_CLK);
    U74HC02 U7040(__A07_NET_195, RT_n, RCH_n, __A07_NET_153, WT_n, WCH_n, GND, WCH_n, CT_n, __A07_NET_151,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1) U7041(__A07_NET_195, __A07_2__RCHG_n, __A07_NET_153, WCHG_n, __A07_NET_151, CCHG_n, GND, __A07_NET_152, WG_n, __A07_1__WGA_n, __A07_NET_152, U2BBKG_n, U2BBK, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8001(__A08_NET_205, A2XG_n, __A08_1___A1_n, __A08_NET_200, WYLOG_n, WL01_n, GND, WL16_n, WYDLOG_n, __A08_NET_199, __A08_1__Y1_n, CUG, __A08_1__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8002(PONEX, __A08_NET_205, __A08_1__X1_n, CLXC, CUG, __A08_1__X1, GND, __A08_1__Y1_n, __A08_NET_200, __A08_NET_199, __A08_1__Y1, __A08_1__X1_n, __A08_1__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8003(__A08_NET_209, __A08_1__X1_n, __A08_1__Y1_n, XUY01_n, __A08_1__X1, __A08_1__Y1, GND, __A08_NET_209, XUY01_n, __A08_NET_207, __A08_NET_209, SUMA01_n, __A08_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8004( ,  , SUMA01_n, SUMB01_n, RULOG_n, __A08_NET_187, GND, __A08_NET_191, __A08_2___XUY1, XUY01_n, CI01_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U8005(CI01_n, __A08_NET_206, G01_n, GEM01, RL01_n, __A08_1___WL1, GND, WL01_n, __A08_1___WL1, __A08_1___MWL1, RL01_n, __A08_NET_157, __A08_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8006(SUMB01_n, __A08_NET_207, __A08_NET_206, __A08_NET_190, WAG_n, WL01_n, GND, WL03_n, WALSG_n, __A08_NET_192, __A08_1___A1_n, CAG, __A08_NET_188, VCC, SIM_RST, SIM_CLK);
    assign __A08_2___CO_IN = __A08_2___CO_IN_U8007_2;
    assign RL01_n = RL01_n_U8007_4;
    assign L01_n = L01_n_U8007_6;
    assign __A08_1___Z1_n = __A08_1___Z1_n_U8007_8;
    assign RL01_n = RL01_n_U8007_10;
    assign RL01_n = RL01_n_U8007_12;
    U74LVC07 U8007(__A08_NET_191, __A08_2___CO_IN_U8007_2, __A08_NET_185, RL01_n_U8007_4, __A08_NET_198, L01_n_U8007_6, GND, __A08_1___Z1_n_U8007_8, __A08_NET_221, RL01_n_U8007_10, __A08_NET_222, RL01_n_U8007_12, __A08_NET_220, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8008(__A08_NET_186, RAG_n, __A08_1___A1_n, __A08_NET_189, WLG_n, WL01_n, GND, __A08_2___G2_n, G2LSG_n, __A08_NET_196, L01_n, CLG1G, __A08_NET_197, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8009( ,  ,  , __A08_NET_194, WQG_n, WL01_n, GND, __A08_NET_194, __A08_NET_193, __A08_1___Q1_n, __A08_1___Q1_n, CQG, __A08_NET_193, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8010(__A08_NET_195, RQG_n, __A08_1___Q1_n, __A08_NET_224, WZG_n, WL01_n, GND, __A08_NET_224, __A08_NET_223, __A08_NET_221, __A08_1___Z1_n, CZG, __A08_NET_223, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8011(__A08_1___RL_OUT_1, __A08_NET_195, MDT01, RB1, R15, __A08_NET_220, GND, __A08_NET_227, __A08_NET_225, __A08_NET_226, __A08_NET_212, __A08_NET_222, __A08_NET_219, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8012(__A08_NET_219, RZG_n, __A08_1___Z1_n, __A08_NET_228, WBG_n, WL01_n, GND, __A08_NET_228, __A08_NET_229, __A08_1___B1_n, __A08_1___B1_n, CBG, __A08_NET_229, VCC, SIM_RST, SIM_CLK);
    assign __A08_2___CO_IN = __A08_2___CO_IN_U8013_2;
    assign RL01_n = RL01_n_U8013_4;
    assign G01_n = G01_n_U8013_6;
    assign G01_n = G01_n_U8013_8;
    assign RL02_n = RL02_n_U8013_10;
    assign L02_n = L02_n_U8013_12;
    U74LVC07 U8013(__A08_NET_170, __A08_2___CO_IN_U8013_2, __A08_NET_227, RL01_n_U8013_4, __A08_NET_211, G01_n_U8013_6, GND, G01_n_U8013_8, __A08_NET_210, RL02_n_U8013_10, __A08_NET_137, L02_n_U8013_12, __A08_NET_147, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8014(__A08_NET_225, RBLG_n, __A08_1___B1_n, __A08_NET_226, __A08_NET_229, RCG_n, GND, WL16_n, WG3G_n, __A08_NET_216, WL02_n, WG4G_n, __A08_NET_215, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8015(__A08_NET_190, __A08_NET_192, __A08_NET_187, __A08_NET_186, CH01, __A08_NET_185, GND, __A08_NET_198, __A08_NET_189, __A08_NET_196, __A08_NET_197, __A08_1___A1_n, __A08_NET_188, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8016(__A08_NET_214, L2GDG_n, MCRO_n, __A08_NET_213, WG1G_n, WL01_n, GND, G01_n, CGG, G01, RGG_n, G01_n, __A08_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U8017(__A08_NET_214, __A08_NET_213, WHOMPA, __A08_2___XUY2, XUY02_n, __A08_NET_170, GND, __A08_1___RL_OUT_1, RLG_n, L01_n, GND, __A08_NET_210, G01, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U8018(__A08_NET_211, G01ED, SA01, __A08_NET_216, __A08_NET_215,  , GND,  , G02ED, SA02, __A08_NET_164, __A08_NET_163, __A08_NET_162, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8019(__A08_NET_158, A2XG_n, __A08_1___A2_n, __A08_NET_160, WYLOG_n, WL02_n, GND, WL01_n, WYDG_n, __A08_NET_159, __A08_1__Y2_n, CUG, __A08_1__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8020(TWOX, __A08_NET_158, __A08_1__X2_n, CLXC, CUG, __A08_1__X2, GND, __A08_1__Y2_n, __A08_NET_160, __A08_NET_159, __A08_1__Y2, __A08_1__X2_n, __A08_1__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8021(__A08_NET_152, __A08_1__X2_n, __A08_1__Y2_n, XUY02_n, __A08_1__X2, __A08_1__Y2, GND,  ,  ,  , __A08_NET_152, XUY02_n, __A08_NET_155, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8022( ,  , __A08_NET_152, SUMA02_n, GND, __A08_2___CI_IN, GND, __A08_NET_156, SUMA02_n, SUMB02_n, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U8023(SUMB02_n, __A08_NET_155, __A08_NET_157, __A08_NET_141, WAG_n, WL02_n, GND, WL04_n, WALSG_n, __A08_NET_140, __A08_1___A2_n, CAG, __A08_NET_139, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8024(__A08_NET_141, __A08_NET_140, __A08_NET_156, __A08_NET_142, CH02, __A08_NET_137, GND, __A08_NET_147, __A08_NET_175, __A08_NET_176, __A08_NET_177, __A08_1___A2_n, __A08_NET_139, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8025(__A08_NET_142, RAG_n, __A08_1___A2_n, __A08_NET_175, WLG_n, WL02_n, GND, G05_n, G2LSG_n, __A08_NET_176, L02_n, CLG1G, __A08_NET_177, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8026(RLG_n, L02_n, __A08_1___RL_OUT_2, __A08_NET_143, __A08_NET_149, __A08_NET_148, GND, __A08_NET_138, MDT02, R1C, RB2, __A08_1___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8027(__A08_NET_179, WQG_n, WL02_n, __A08_1___Q2_n, __A08_NET_179, __A08_NET_178, GND, __A08_1___Q2_n, CQG, __A08_NET_178, RQG_n, __A08_1___Q2_n, __A08_NET_143, VCC, SIM_RST, SIM_CLK);
    assign RL02_n = RL02_n_U8028_2;
    assign __A08_1___Z2_n = __A08_1___Z2_n_U8028_4;
    assign RL02_n = RL02_n_U8028_6;
    assign RL02_n = RL02_n_U8028_8;
    assign __A08_1___G2_n = __A08_1___G2_n_U8028_10;
    assign __A08_1___G2_n = __A08_1___G2_n_U8028_12;
    U74LVC07 U8028(__A08_NET_148, RL02_n_U8028_2, __A08_NET_145, __A08_1___Z2_n_U8028_4, __A08_NET_138, RL02_n_U8028_6, GND, RL02_n_U8028_8, __A08_NET_180, __A08_1___G2_n_U8028_10, __A08_NET_162, __A08_1___G2_n_U8028_12, __A08_NET_169, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8029(__A08_NET_144, WZG_n, WL02_n, __A08_NET_145, __A08_NET_144, __A08_NET_146, GND, __A08_1___Z2_n, CZG, __A08_NET_146, RZG_n, __A08_1___Z2_n, __A08_NET_149, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8030(__A08_NET_183, WBG_n, WL02_n, __A08_1___B2_n, __A08_NET_183, __A08_NET_184, GND, __A08_1___B2_n, CBG, __A08_NET_184, RBLG_n, __A08_1___B2_n, __A08_NET_182, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U8031(__A08_NET_182, __A08_NET_181, __A08_NET_168, __A08_NET_167, G02, __A08_NET_169, GND, __A08_NET_263, GND, XUY06_n, __A08_2___XUY2, __A08_NET_180, __A08_NET_161, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8032(__A08_NET_181, __A08_NET_184, RCG_n, __A08_NET_164, WL01_n, WG3G_n, GND, WL03_n, WG4G_n, __A08_NET_163, L2GDG_n, L01_n, __A08_NET_168, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8033(__A08_NET_167, WG1G_n, WL02_n, G02, __A08_1___G2_n, CGG, GND, RGG_n, __A08_1___G2_n, __A08_NET_161,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U8034(__A08_1___G2_n, GEM02, RL02_n, __A08_1___WL2, __A08_1___WL2, WL02_n, GND, __A08_1___MWL2, RL02_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U8035(__A08_NET_298, A2XG_n, __A08_2___A1_n, __A08_NET_294, WYLOG_n, WL03_n, GND, WL02_n, WYDG_n, __A08_NET_293, __A08_2__Y1_n, CUG, __A08_2__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8036(MONEX, __A08_NET_298, __A08_2__X1_n, CLXC, CUG, __A08_2__X1, GND, __A08_2__Y1_n, __A08_NET_294, __A08_NET_293, __A08_2__Y1, __A08_2__X1_n, __A08_2__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8037(__A08_NET_302, __A08_2__X1_n, __A08_2__Y1_n, __A08_2___XUY1, __A08_2__X1, __A08_2__Y1, GND, __A08_NET_302, __A08_2___XUY1, __A08_NET_299, __A08_NET_302, SUMA03_n, __A08_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8038( ,  , SUMA03_n, SUMB03_n, RULOG_n, __A08_NET_280, GND, __A08_NET_284, XUY05_n, __A08_2___XUY1, __A08_2___CI_IN,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U8039(__A08_2___CI_IN, __A08_NET_300, __A08_2___G1_n, GEM03, RL03_n, __A08_2___WL1, GND, WL03_n, __A08_2___WL1, __A08_2___MWL1, RL03_n, __A08_NET_250, __A08_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8040(SUMB03_n, __A08_NET_299, __A08_NET_300, __A08_NET_283, WAG_n, WL03_n, GND, WL05_n, WALSG_n, __A08_NET_285, __A08_2___A1_n, CAG, __A08_NET_281, VCC, SIM_RST, SIM_CLK);
    assign CO06 = CO06_U8041_2;
    assign RL03_n = RL03_n_U8041_4;
    assign __A08_2___L1_n = __A08_2___L1_n_U8041_6;
    assign __A08_2___Z1_n = __A08_2___Z1_n_U8041_8;
    assign RL03_n = RL03_n_U8041_10;
    assign RL03_n = RL03_n_U8041_12;
    U74LVC07 U8041(__A08_NET_284, CO06_U8041_2, __A08_NET_279, RL03_n_U8041_4, __A08_NET_291, __A08_2___L1_n_U8041_6, GND, __A08_2___Z1_n_U8041_8, __A08_NET_314, RL03_n_U8041_10, __A08_NET_315, RL03_n_U8041_12, __A08_NET_313, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8042(__A08_NET_283, __A08_NET_285, __A08_NET_280, __A08_NET_278, CH03, __A08_NET_279, GND, __A08_NET_291, __A08_NET_282, __A08_NET_289, __A08_NET_290, __A08_2___A1_n, __A08_NET_281, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8043(__A08_NET_278, RAG_n, __A08_2___A1_n, __A08_NET_282, WLG_n, WL03_n, GND, G06_n, G2LSG_n, __A08_NET_289, __A08_2___L1_n, CLG1G, __A08_NET_290, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8044( ,  ,  ,  ,  ,  , GND, __A08_2___RL_OUT_1, RLG_n, __A08_2___L1_n, GND,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8045( ,  ,  , __A08_NET_287, WQG_n, WL03_n, GND, __A08_NET_287, __A08_NET_286, __A08_2___Q1_n, __A08_2___Q1_n, CQG, __A08_NET_286, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8046(__A08_NET_288, RQG_n, __A08_2___Q1_n, __A08_NET_317, WZG_n, WL03_n, GND, __A08_NET_317, __A08_NET_316, __A08_NET_314, __A08_2___Z1_n, CZG, __A08_NET_316, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8047(__A08_NET_312, RZG_n, __A08_2___Z1_n, __A08_NET_321, WBG_n, WL03_n, GND, __A08_NET_321, __A08_NET_322, __A08_2___B1_n, __A08_2___B1_n, CBG, __A08_NET_322, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8048(__A08_NET_319, RBLG_n, __A08_2___B1_n, __A08_NET_320, __A08_NET_322, RCG_n, GND, WL02_n, WG3G_n, __A08_NET_309, WL04_n, WG4G_n, __A08_NET_308, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8049(__A08_2___RL_OUT_1, __A08_NET_288, MDT03, R1C, R15, __A08_NET_313, GND, __A08_NET_318, __A08_NET_319, __A08_NET_320, __A08_NET_305, __A08_NET_315, __A08_NET_312, VCC, SIM_RST, SIM_CLK);
    assign CO06 = CO06_U8050_2;
    assign RL03_n = RL03_n_U8050_4;
    assign __A08_2___G1_n = __A08_2___G1_n_U8050_6;
    assign __A08_2___G1_n = __A08_2___G1_n_U8050_8;
    assign RL04_n = RL04_n_U8050_10;
    assign L04_n = L04_n_U8050_12;
    U74LVC07 U8050(__A08_NET_263, CO06_U8050_2, __A08_NET_318, RL03_n_U8050_4, __A08_NET_304, __A08_2___G1_n_U8050_6, GND, __A08_2___G1_n_U8050_8, __A08_NET_303, RL04_n_U8050_10, __A08_NET_230, L04_n_U8050_12, __A08_NET_240, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8051(__A08_NET_307, L2GDG_n, L02_n, __A08_NET_306, WG1G_n, WL03_n, GND, __A08_2___G1_n, CGG, G03, RGG_n, __A08_2___G1_n, __A08_NET_305, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U8052(__A08_NET_304, G03ED, SA03, __A08_NET_309, __A08_NET_308,  , GND,  , G04ED, SA04, __A08_NET_257, __A08_NET_256, __A08_NET_255, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U8053(__A08_NET_307, __A08_NET_306,  ,  ,  ,  , GND,  ,  ,  ,  , __A08_NET_303, G03, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8054(__A08_NET_251, A2XG_n, __A08_2___A2_n, __A08_NET_253, WYLOG_n, WL04_n, GND, WL03_n, WYDG_n, __A08_NET_252, __A08_2__Y2_n, CUG, __A08_2__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8055(MONEX, __A08_NET_251, __A08_2__X2_n, CLXC, CUG, __A08_2__X2, GND, __A08_2__Y2_n, __A08_NET_253, __A08_NET_252, __A08_2__Y2, __A08_2__X2_n, __A08_2__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8056(__A08_NET_245, __A08_2__X2_n, __A08_2__Y2_n, __A08_2___XUY2, __A08_2__X2, __A08_2__Y2, GND,  ,  ,  , __A08_NET_245, __A08_2___XUY2, __A08_NET_248, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8057( ,  , __A08_NET_245, __A08_2___SUMA2, __A08_2___CO_IN, CI05_n, GND, __A08_NET_249, __A08_2___SUMA2, __A08_2___SUMB2, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U8058(__A08_2___SUMB2, __A08_NET_248, __A08_NET_250, __A08_NET_234, WAG_n, WL04_n, GND, WL06_n, WALSG_n, __A08_NET_233, __A08_2___A2_n, CAG, __A08_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8059(__A08_NET_234, __A08_NET_233, __A08_NET_249, __A08_NET_235, CH04, __A08_NET_230, GND, __A08_NET_240, __A08_NET_268, __A08_NET_269, __A08_NET_270, __A08_2___A2_n, __A08_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8060(__A08_NET_235, RAG_n, __A08_2___A2_n, __A08_NET_268, WLG_n, WL04_n, GND, G07_n, G2LSG_n, __A08_NET_269, L04_n, CLG1G, __A08_NET_270, VCC, SIM_RST, SIM_CLK);
    U74HC27 U8061(RLG_n, L04_n, __A08_2___RL_OUT_2, __A08_NET_236, __A08_NET_242, __A08_NET_241, GND, __A08_NET_231, MDT04, R1C, R15, __A08_2___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8062(__A08_NET_272, WQG_n, WL04_n, __A08_2___Q2_n, __A08_NET_272, __A08_NET_271, GND, __A08_2___Q2_n, CQG, __A08_NET_271, RQG_n, __A08_2___Q2_n, __A08_NET_236, VCC, SIM_RST, SIM_CLK);
    assign RL04_n = RL04_n_U8063_2;
    assign __A08_2___Z2_n = __A08_2___Z2_n_U8063_4;
    assign RL04_n = RL04_n_U8063_6;
    assign RL04_n = RL04_n_U8063_8;
    assign __A08_2___G2_n = __A08_2___G2_n_U8063_10;
    assign __A08_2___G2_n = __A08_2___G2_n_U8063_12;
    U74LVC07 U8063(__A08_NET_241, RL04_n_U8063_2, __A08_NET_238, __A08_2___Z2_n_U8063_4, __A08_NET_231, RL04_n_U8063_6, GND, RL04_n_U8063_8, __A08_NET_273, __A08_2___G2_n_U8063_10, __A08_NET_255, __A08_2___G2_n_U8063_12, __A08_NET_262, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8064(__A08_NET_237, WZG_n, WL04_n, __A08_NET_238, __A08_NET_237, __A08_NET_239, GND, __A08_2___Z2_n, CZG, __A08_NET_239, RZG_n, __A08_2___Z2_n, __A08_NET_242, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8065(__A08_NET_276, WBG_n, WL04_n, __A08_2___B2_n, __A08_NET_276, __A08_NET_277, GND, __A08_2___B2_n, CBG, __A08_NET_277, RBLG_n, __A08_2___B2_n, __A08_NET_275, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U8066(__A08_NET_275, __A08_NET_274, __A08_NET_261, __A08_NET_260, G04, __A08_NET_262, GND,  ,  ,  ,  , __A08_NET_273, __A08_NET_254, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8067(__A08_NET_274, __A08_NET_277, RCG_n, __A08_NET_257, WL03_n, WG3G_n, GND, WL05_n, WG4G_n, __A08_NET_256, L2GDG_n, __A08_2___L1_n, __A08_NET_261, VCC, SIM_RST, SIM_CLK);
    U74HC02 U8068(__A08_NET_260, WG1G_n, WL04_n, G04, __A08_2___G2_n, CGG, GND, RGG_n, __A08_2___G2_n, __A08_NET_254,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U8069(__A08_2___G2_n, GEM04, RL04_n, __A08_2___WL2, __A08_2___WL2, WL04_n, GND, __A08_2___MWL2, RL04_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC4002 U8070(SUMA01_n, __A08_NET_209, XUY01_n, CI01_n, GND,  , GND,  , __A08_NET_152, XUY02_n, __A08_1___CI_INTERNAL, WHOMP, SUMA02_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U8071(SUMA03_n, __A08_NET_302, __A08_2___XUY1, __A08_2___CI_IN, GND,  , GND,  , __A08_NET_245, __A08_2___XUY2, __A08_2___CI_INTERNAL, WHOMP, __A08_2___SUMA2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9001(__A09_NET_198, A2XG_n, __A09_1___A1_n, __A09_NET_193, WYLOG_n, WL05_n, GND, WL04_n, WYDG_n, __A09_NET_192, __A09_1__Y1_n, CUG, __A09_1__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9002(MONEX, __A09_NET_198, __A09_1__X1_n, CLXC, CUG, __A09_1__X1, GND, __A09_1__Y1_n, __A09_NET_193, __A09_NET_192, __A09_1__Y1, __A09_1__X1_n, __A09_1__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9003(__A09_NET_202, __A09_1__X1_n, __A09_1__Y1_n, XUY05_n, __A09_1__X1, __A09_1__Y1, GND, __A09_NET_202, XUY05_n, __A09_NET_200, __A09_NET_202, __A09_1___SUMA1, __A09_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9004( ,  , __A09_1___SUMA1, __A09_1___SUMB1, RULOG_n, __A09_NET_180, GND, __A09_NET_184, __A09_2___XUY1, XUY05_n, CI05_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U9005(CI05_n, __A09_NET_199, G05_n, GEM05, RL05_n, __A09_1___WL1, GND, WL05_n, __A09_1___WL1, __A09_1___MWL1, RL05_n, __A09_NET_150, __A09_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9006(__A09_1___SUMB1, __A09_NET_200, __A09_NET_199, __A09_NET_183, WAG_n, WL05_n, GND, WL07_n, WALSG_n, __A09_NET_185, __A09_1___A1_n, CAG, __A09_NET_181, VCC, SIM_RST, SIM_CLK);
    assign __A09_2___CO_IN = __A09_2___CO_IN_U9007_2;
    assign RL05_n = RL05_n_U9007_4;
    assign __A09_1___L1_n = __A09_1___L1_n_U9007_6;
    assign __A09_1___Z1_n = __A09_1___Z1_n_U9007_8;
    assign RL05_n = RL05_n_U9007_10;
    assign RL05_n = RL05_n_U9007_12;
    U74LVC07 U9007(__A09_NET_184, __A09_2___CO_IN_U9007_2, __A09_NET_178, RL05_n_U9007_4, __A09_NET_191, __A09_1___L1_n_U9007_6, GND, __A09_1___Z1_n_U9007_8, __A09_NET_214, RL05_n_U9007_10, __A09_NET_215, RL05_n_U9007_12, __A09_NET_213, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9008(__A09_NET_179, RAG_n, __A09_1___A1_n, __A09_NET_182, WLG_n, WL05_n, GND, __A09_2___G2_n, G2LSG_n, __A09_NET_189, __A09_1___L1_n, CLG1G, __A09_NET_190, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9009( ,  ,  , __A09_NET_187, WQG_n, WL05_n, GND, __A09_NET_187, __A09_NET_186, __A09_1___Q1_n, __A09_1___Q1_n, CQG, __A09_NET_186, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9010(__A09_NET_188, RQG_n, __A09_1___Q1_n, __A09_NET_217, WZG_n, WL05_n, GND, __A09_NET_217, __A09_NET_216, __A09_NET_214, __A09_1___Z1_n, CZG, __A09_NET_216, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9011(__A09_1___RL_OUT_1, __A09_NET_188, MDT05, R1C, GND, __A09_NET_213, GND, __A09_NET_220, __A09_NET_218, __A09_NET_219, __A09_NET_205, __A09_NET_215, __A09_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9012(__A09_NET_212, RZG_n, __A09_1___Z1_n, __A09_NET_221, WBG_n, WL05_n, GND, __A09_NET_221, __A09_NET_222, __A09_1___B1_n, __A09_1___B1_n, CBG, __A09_NET_222, VCC, SIM_RST, SIM_CLK);
    assign __A09_2___CO_IN = __A09_2___CO_IN_U9013_2;
    assign RL05_n = RL05_n_U9013_4;
    assign G05_n = G05_n_U9013_6;
    assign G05_n = G05_n_U9013_8;
    assign RL06_n = RL06_n_U9013_10;
    assign __A09_1___L2_n = __A09_1___L2_n_U9013_12;
    U74LVC07 U9013(__A09_NET_163, __A09_2___CO_IN_U9013_2, __A09_NET_220, RL05_n_U9013_4, __A09_NET_204, G05_n_U9013_6, GND, G05_n_U9013_8, __A09_NET_203, RL06_n_U9013_10, __A09_NET_130, __A09_1___L2_n_U9013_12, __A09_NET_140, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9014(__A09_NET_218, RBLG_n, __A09_1___B1_n, __A09_NET_219, __A09_NET_222, RCG_n, GND, WL04_n, WG3G_n, __A09_NET_209, WL06_n, WG4G_n, __A09_NET_208, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9015(__A09_NET_183, __A09_NET_185, __A09_NET_180, __A09_NET_179, CH05, __A09_NET_178, GND, __A09_NET_191, __A09_NET_182, __A09_NET_189, __A09_NET_190, __A09_1___A1_n, __A09_NET_181, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9016(__A09_NET_207, L2GDG_n, L04_n, __A09_NET_206, WG1G_n, WL05_n, GND, G05_n, CGG, G05, RGG_n, G05_n, __A09_NET_205, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U9017(__A09_NET_207, __A09_NET_206, GND, __A09_2___XUY2, XUY06_n, __A09_NET_163, GND, __A09_1___RL_OUT_1, RLG_n, __A09_1___L1_n, GND, __A09_NET_203, G05, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U9018(__A09_NET_204, G05ED, SA05, __A09_NET_209, __A09_NET_208,  , GND,  , G06ED, SA06, __A09_NET_157, __A09_NET_156, __A09_NET_155, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9019(__A09_NET_151, A2XG_n, __A09_1___A2_n, __A09_NET_153, WYLOG_n, WL06_n, GND, WL05_n, WYDG_n, __A09_NET_152, __A09_1__Y2_n, CUG, __A09_1__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9020(MONEX, __A09_NET_151, __A09_1__X2_n, CLXC, CUG, __A09_1__X2, GND, __A09_1__Y2_n, __A09_NET_153, __A09_NET_152, __A09_1__Y2, __A09_1__X2_n, __A09_1__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9021(__A09_NET_145, __A09_1__X2_n, __A09_1__Y2_n, XUY06_n, __A09_1__X2, __A09_1__Y2, GND,  ,  ,  , __A09_NET_145, XUY06_n, __A09_NET_148, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9022( ,  , __A09_NET_145, __A09_1___SUMA2, CO06, __A09_2___CI_IN, GND, __A09_NET_149, __A09_1___SUMA2, __A09_1___SUMB2, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U9023(__A09_1___SUMB2, __A09_NET_148, __A09_NET_150, __A09_NET_134, WAG_n, WL06_n, GND, WL08_n, WALSG_n, __A09_NET_133, __A09_1___A2_n, CAG, __A09_NET_132, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9024(__A09_NET_134, __A09_NET_133, __A09_NET_149, __A09_NET_135, CH06, __A09_NET_130, GND, __A09_NET_140, __A09_NET_168, __A09_NET_169, __A09_NET_170, __A09_1___A2_n, __A09_NET_132, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9025(__A09_NET_135, RAG_n, __A09_1___A2_n, __A09_NET_168, WLG_n, WL06_n, GND, G09_n, G2LSG_n, __A09_NET_169, __A09_1___L2_n, CLG1G, __A09_NET_170, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9026(RLG_n, __A09_1___L2_n, __A09_1___RL_OUT_2, __A09_NET_136, __A09_NET_142, __A09_NET_141, GND, __A09_NET_131, MDT06, R1C, GND, __A09_1___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9027(__A09_NET_172, WQG_n, WL06_n, __A09_1___Q2_n, __A09_NET_172, __A09_NET_171, GND, __A09_1___Q2_n, CQG, __A09_NET_171, RQG_n, __A09_1___Q2_n, __A09_NET_136, VCC, SIM_RST, SIM_CLK);
    assign RL06_n = RL06_n_U9028_2;
    assign __A09_1___Z2_n = __A09_1___Z2_n_U9028_4;
    assign RL06_n = RL06_n_U9028_6;
    assign RL06_n = RL06_n_U9028_8;
    assign G06_n = G06_n_U9028_10;
    assign G06_n = G06_n_U9028_12;
    U74LVC07 U9028(__A09_NET_141, RL06_n_U9028_2, __A09_NET_138, __A09_1___Z2_n_U9028_4, __A09_NET_131, RL06_n_U9028_6, GND, RL06_n_U9028_8, __A09_NET_173, G06_n_U9028_10, __A09_NET_155, G06_n_U9028_12, __A09_NET_162, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9029(__A09_NET_137, WZG_n, WL06_n, __A09_NET_138, __A09_NET_137, __A09_NET_139, GND, __A09_1___Z2_n, CZG, __A09_NET_139, RZG_n, __A09_1___Z2_n, __A09_NET_142, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9030(__A09_NET_176, WBG_n, WL06_n, __A09_1___B2_n, __A09_NET_176, __A09_NET_177, GND, __A09_1___B2_n, CBG, __A09_NET_177, RBLG_n, __A09_1___B2_n, __A09_NET_175, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U9031(__A09_NET_175, __A09_NET_174, __A09_NET_161, __A09_NET_160, G06, __A09_NET_162, GND, __A09_NET_256, GND, XUY10_n, __A09_2___XUY2, __A09_NET_173, __A09_NET_154, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9032(__A09_NET_174, __A09_NET_177, RCG_n, __A09_NET_157, WL05_n, WG3G_n, GND, WL07_n, WG4G_n, __A09_NET_156, L2GDG_n, __A09_1___L1_n, __A09_NET_161, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9033(__A09_NET_160, WG1G_n, WL06_n, G06, G06_n, CGG, GND, RGG_n, G06_n, __A09_NET_154,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U9034(G06_n, GEM06, RL06_n, __A09_1___WL2, __A09_1___WL2, WL06_n, GND, __A09_1___MWL2, RL06_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U9035(__A09_NET_291, A2XG_n, __A09_2___A1_n, __A09_NET_287, WYLOG_n, WL07_n, GND, WL06_n, WYDG_n, __A09_NET_286, __A09_2__Y1_n, CUG, __A09_2__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9036(MONEX, __A09_NET_291, __A09_2__X1_n, CLXC, CUG, __A09_2__X1, GND, __A09_2__Y1_n, __A09_NET_287, __A09_NET_286, __A09_2__Y1, __A09_2__X1_n, __A09_2__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9037(__A09_NET_295, __A09_2__X1_n, __A09_2__Y1_n, __A09_2___XUY1, __A09_2__X1, __A09_2__Y1, GND, __A09_NET_295, __A09_2___XUY1, __A09_NET_292, __A09_NET_295, __A09_2___SUMA1, __A09_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9038( ,  , __A09_2___SUMA1, __A09_2___SUMB1, RULOG_n, __A09_NET_273, GND, __A09_NET_277, XUY09_n, __A09_2___XUY1, __A09_2___CI_IN,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U9039(__A09_2___CI_IN, __A09_NET_293, G07_n, GEM07, __A09_2___RL1_n, __A09_2___WL1, GND, WL07_n, __A09_2___WL1, __A09_2___MWL1, __A09_2___RL1_n, __A09_NET_243, __A09_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9040(__A09_2___SUMB1, __A09_NET_292, __A09_NET_293, __A09_NET_276, WAG_n, WL07_n, GND, WL09_n, WALSG_n, __A09_NET_278, __A09_2___A1_n, CAG, __A09_NET_274, VCC, SIM_RST, SIM_CLK);
    assign CO10 = CO10_U9041_2;
    assign __A09_2___RL1_n = __A09_2___RL1_n_U9041_4;
    assign __A09_2___L1_n = __A09_2___L1_n_U9041_6;
    assign __A09_2___Z1_n = __A09_2___Z1_n_U9041_8;
    assign __A09_2___RL1_n = __A09_2___RL1_n_U9041_10;
    assign __A09_2___RL1_n = __A09_2___RL1_n_U9041_12;
    U74LVC07 U9041(__A09_NET_277, CO10_U9041_2, __A09_NET_272, __A09_2___RL1_n_U9041_4, __A09_NET_284, __A09_2___L1_n_U9041_6, GND, __A09_2___Z1_n_U9041_8, __A09_NET_307, __A09_2___RL1_n_U9041_10, __A09_NET_308, __A09_2___RL1_n_U9041_12, __A09_NET_306, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9042(__A09_NET_276, __A09_NET_278, __A09_NET_273, __A09_NET_271, CH07, __A09_NET_272, GND, __A09_NET_284, __A09_NET_275, __A09_NET_282, __A09_NET_283, __A09_2___A1_n, __A09_NET_274, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9043(__A09_NET_271, RAG_n, __A09_2___A1_n, __A09_NET_275, WLG_n, WL07_n, GND, G10_n, G2LSG_n, __A09_NET_282, __A09_2___L1_n, CLG1G, __A09_NET_283, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9044( ,  ,  ,  ,  ,  , GND, __A09_2___RL_OUT_1, RLG_n, __A09_2___L1_n, GND,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9045( ,  ,  , __A09_NET_280, WQG_n, WL07_n, GND, __A09_NET_280, __A09_NET_279, __A09_2___Q1_n, __A09_2___Q1_n, CQG, __A09_NET_279, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9046(__A09_NET_281, RQG_n, __A09_2___Q1_n, __A09_NET_310, WZG_n, WL07_n, GND, __A09_NET_310, __A09_NET_309, __A09_NET_307, __A09_2___Z1_n, CZG, __A09_NET_309, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9047(__A09_NET_305, RZG_n, __A09_2___Z1_n, __A09_NET_314, WBG_n, WL07_n, GND, __A09_NET_314, __A09_NET_315, __A09_2___B1_n, __A09_2___B1_n, CBG, __A09_NET_315, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9048(__A09_NET_312, RBLG_n, __A09_2___B1_n, __A09_NET_313, __A09_NET_315, RCG_n, GND, WL06_n, WG3G_n, __A09_NET_302, WL08_n, WG4G_n, __A09_NET_301, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9049(__A09_2___RL_OUT_1, __A09_NET_281, MDT07, R1C, GND, __A09_NET_306, GND, __A09_NET_311, __A09_NET_312, __A09_NET_313, __A09_NET_298, __A09_NET_308, __A09_NET_305, VCC, SIM_RST, SIM_CLK);
    assign CO10 = CO10_U9050_2;
    assign __A09_2___RL1_n = __A09_2___RL1_n_U9050_4;
    assign G07_n = G07_n_U9050_6;
    assign G07_n = G07_n_U9050_8;
    assign __A09_2___RL2_n = __A09_2___RL2_n_U9050_10;
    assign L08_n = L08_n_U9050_12;
    U74LVC07 U9050(__A09_NET_256, CO10_U9050_2, __A09_NET_311, __A09_2___RL1_n_U9050_4, __A09_NET_297, G07_n_U9050_6, GND, G07_n_U9050_8, __A09_NET_296, __A09_2___RL2_n_U9050_10, __A09_NET_223, L08_n_U9050_12, __A09_NET_233, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9051(__A09_NET_300, L2GDG_n, __A09_1___L2_n, __A09_NET_299, WG1G_n, WL07_n, GND, G07_n, CGG, G07, RGG_n, G07_n, __A09_NET_298, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U9052(__A09_NET_297, G07ED, SA07, __A09_NET_302, __A09_NET_301,  , GND,  , GND, SA08, __A09_NET_250, __A09_NET_249, __A09_NET_248, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U9053(__A09_NET_300, __A09_NET_299,  ,  ,  ,  , GND,  ,  ,  ,  , __A09_NET_296, G07, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9054(__A09_NET_244, A2XG_n, __A09_2___A2_n, __A09_NET_246, WYLOG_n, WL08_n, GND, WL07_n, WYDG_n, __A09_NET_245, __A09_2__Y2_n, CUG, __A09_2__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9055(MONEX, __A09_NET_244, __A09_2__X2_n, CLXC, CUG, __A09_2__X2, GND, __A09_2__Y2_n, __A09_NET_246, __A09_NET_245, __A09_2__Y2, __A09_2__X2_n, __A09_2__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9056(__A09_NET_238, __A09_2__X2_n, __A09_2__Y2_n, __A09_2___XUY2, __A09_2__X2, __A09_2__Y2, GND,  ,  ,  , __A09_NET_238, __A09_2___XUY2, __A09_NET_241, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9057( ,  , __A09_NET_238, __A09_2___SUMA2, __A09_2___CO_IN, CI09_n, GND, __A09_NET_242, __A09_2___SUMA2, __A09_2___SUMB2, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U9058(__A09_2___SUMB2, __A09_NET_241, __A09_NET_243, __A09_NET_227, WAG_n, WL08_n, GND, WL10_n, WALSG_n, __A09_NET_226, __A09_2___A2_n, CAG, __A09_NET_225, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9059(__A09_NET_227, __A09_NET_226, __A09_NET_242, __A09_NET_228, CH08, __A09_NET_223, GND, __A09_NET_233, __A09_NET_261, __A09_NET_262, __A09_NET_263, __A09_2___A2_n, __A09_NET_225, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9060(__A09_NET_228, RAG_n, __A09_2___A2_n, __A09_NET_261, WLG_n, WL08_n, GND, G11_n, G2LSG_n, __A09_NET_262, L08_n, CLG1G, __A09_NET_263, VCC, SIM_RST, SIM_CLK);
    U74HC27 U9061(RLG_n, L08_n, __A09_2___RL_OUT_2, __A09_NET_229, __A09_NET_235, __A09_NET_234, GND, __A09_NET_224, MDT08, R1C, GND, __A09_2___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9062(__A09_NET_265, WQG_n, WL08_n, __A09_2___Q2_n, __A09_NET_265, __A09_NET_264, GND, __A09_2___Q2_n, CQG, __A09_NET_264, RQG_n, __A09_2___Q2_n, __A09_NET_229, VCC, SIM_RST, SIM_CLK);
    assign __A09_2___RL2_n = __A09_2___RL2_n_U9063_2;
    assign __A09_2___Z2_n = __A09_2___Z2_n_U9063_4;
    assign __A09_2___RL2_n = __A09_2___RL2_n_U9063_6;
    assign __A09_2___RL2_n = __A09_2___RL2_n_U9063_8;
    assign __A09_2___G2_n = __A09_2___G2_n_U9063_10;
    assign __A09_2___G2_n = __A09_2___G2_n_U9063_12;
    U74LVC07 U9063(__A09_NET_234, __A09_2___RL2_n_U9063_2, __A09_NET_231, __A09_2___Z2_n_U9063_4, __A09_NET_224, __A09_2___RL2_n_U9063_6, GND, __A09_2___RL2_n_U9063_8, __A09_NET_266, __A09_2___G2_n_U9063_10, __A09_NET_248, __A09_2___G2_n_U9063_12, __A09_NET_255, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9064(__A09_NET_230, WZG_n, WL08_n, __A09_NET_231, __A09_NET_230, __A09_NET_232, GND, __A09_2___Z2_n, CZG, __A09_NET_232, RZG_n, __A09_2___Z2_n, __A09_NET_235, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9065(__A09_NET_269, WBG_n, WL08_n, __A09_2___B2_n, __A09_NET_269, __A09_NET_270, GND, __A09_2___B2_n, CBG, __A09_NET_270, RBLG_n, __A09_2___B2_n, __A09_NET_268, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U9066(__A09_NET_268, __A09_NET_267, __A09_NET_254, __A09_NET_253, G08, __A09_NET_255, GND,  ,  ,  ,  , __A09_NET_266, __A09_NET_247, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9067(__A09_NET_267, __A09_NET_270, RCG_n, __A09_NET_250, WL07_n, WG3G_n, GND, WL09_n, WG4G_n, __A09_NET_249, L2GDG_n, __A09_2___L1_n, __A09_NET_254, VCC, SIM_RST, SIM_CLK);
    U74HC02 U9068(__A09_NET_253, WG1G_n, WL08_n, G08, __A09_2___G2_n, CGG, GND, RGG_n, __A09_2___G2_n, __A09_NET_247,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U9069(__A09_2___G2_n, GEM08, __A09_2___RL2_n, __A09_2___WL2, __A09_2___WL2, WL08_n, GND, __A09_2___MWL2, __A09_2___RL2_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC4002 U9070(__A09_1___SUMA1, __A09_NET_202, XUY05_n, CI05_n, GND,  , GND,  , __A09_NET_145, XUY06_n, __A09_1___CI_INTERNAL, GND, __A09_1___SUMA2, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U9071(__A09_2___SUMA1, __A09_NET_295, __A09_2___XUY1, __A09_2___CI_IN, WHOMP,  , GND,  , __A09_NET_238, __A09_2___XUY2, __A09_2___CI_INTERNAL, GND, __A09_2___SUMA2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10001(__A10_NET_197, A2XG_n, __A10_1___A1_n, __A10_NET_192, WYLOG_n, WL09_n, GND, WL08_n, WYDG_n, __A10_NET_191, __A10_1__Y1_n, CUG, __A10_1__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10002(MONEX, __A10_NET_197, __A10_1__X1_n, CLXC, CUG, __A10_1__X1, GND, __A10_1__Y1_n, __A10_NET_192, __A10_NET_191, __A10_1__Y1, __A10_1__X1_n, __A10_1__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10003(__A10_NET_201, __A10_1__X1_n, __A10_1__Y1_n, XUY09_n, __A10_1__X1, __A10_1__Y1, GND, __A10_NET_201, XUY09_n, __A10_NET_199, __A10_NET_201, __A10_1___SUMA1, __A10_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10004( ,  , __A10_1___SUMA1, __A10_1___SUMB1, RULOG_n, __A10_NET_179, GND, __A10_NET_183, __A10_2___XUY1, XUY09_n, CI09_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U10005(CI09_n, __A10_NET_198, G09_n, GEM09, RL09_n, __A10_1___WL1, GND, WL09_n, __A10_1___WL1, __A10_1___MWL1, RL09_n, __A10_NET_149, __A10_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10006(__A10_1___SUMB1, __A10_NET_199, __A10_NET_198, __A10_NET_182, WAG_n, WL09_n, GND, WL11_n, WALSG_n, __A10_NET_184, __A10_1___A1_n, CAG, __A10_NET_180, VCC, SIM_RST, SIM_CLK);
    assign __A10_2___CO_IN = __A10_2___CO_IN_U10007_2;
    assign RL09_n = RL09_n_U10007_4;
    assign __A10_1___L1_n = __A10_1___L1_n_U10007_6;
    assign __A10_1___Z1_n = __A10_1___Z1_n_U10007_8;
    assign RL09_n = RL09_n_U10007_10;
    assign RL09_n = RL09_n_U10007_12;
    U74LVC07 U10007(__A10_NET_183, __A10_2___CO_IN_U10007_2, __A10_NET_177, RL09_n_U10007_4, __A10_NET_190, __A10_1___L1_n_U10007_6, GND, __A10_1___Z1_n_U10007_8, __A10_NET_213, RL09_n_U10007_10, __A10_NET_214, RL09_n_U10007_12, __A10_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10008(__A10_NET_178, RAG_n, __A10_1___A1_n, __A10_NET_181, WLG_n, WL09_n, GND, __A10_2___G2_n, G2LSG_n, __A10_NET_188, __A10_1___L1_n, CLG1G, __A10_NET_189, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U10009( ,  ,  , __A10_NET_186, WQG_n, WL09_n, GND, __A10_NET_186, __A10_NET_185, __A10_1___Q1_n, __A10_1___Q1_n, CQG, __A10_NET_185, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U10010(__A10_NET_187, RQG_n, __A10_1___Q1_n, __A10_NET_216, WZG_n, WL09_n, GND, __A10_NET_216, __A10_NET_215, __A10_NET_213, __A10_1___Z1_n, CZG, __A10_NET_215, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10011(__A10_1___RL_OUT_1, __A10_NET_187, MDT09, R1C, GND, __A10_NET_212, GND, __A10_NET_219, __A10_NET_217, __A10_NET_218, __A10_NET_204, __A10_NET_214, __A10_NET_211, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U10012(__A10_NET_211, RZG_n, __A10_1___Z1_n, __A10_NET_220, WBG_n, WL09_n, GND, __A10_NET_220, __A10_NET_221, __A10_1___B1_n, __A10_1___B1_n, CBG, __A10_NET_221, VCC, SIM_RST, SIM_CLK);
    assign __A10_2___CO_IN = __A10_2___CO_IN_U10013_2;
    assign RL09_n = RL09_n_U10013_4;
    assign G09_n = G09_n_U10013_6;
    assign G09_n = G09_n_U10013_8;
    assign RL10_n = RL10_n_U10013_10;
    assign __A10_1___L2_n = __A10_1___L2_n_U10013_12;
    U74LVC07 U10013(__A10_NET_162, __A10_2___CO_IN_U10013_2, __A10_NET_219, RL09_n_U10013_4, __A10_NET_203, G09_n_U10013_6, GND, G09_n_U10013_8, __A10_NET_202, RL10_n_U10013_10, __A10_NET_129, __A10_1___L2_n_U10013_12, __A10_NET_139, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10014(__A10_NET_217, RBLG_n, __A10_1___B1_n, __A10_NET_218, __A10_NET_221, RCG_n, GND, WL08_n, WG3G_n, __A10_NET_208, WL10_n, WG4G_n, __A10_NET_207, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10015(__A10_NET_182, __A10_NET_184, __A10_NET_179, __A10_NET_178, CH09, __A10_NET_177, GND, __A10_NET_190, __A10_NET_181, __A10_NET_188, __A10_NET_189, __A10_1___A1_n, __A10_NET_180, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10016(__A10_NET_206, L2GDG_n, L08_n, __A10_NET_205, WG1G_n, WL09_n, GND, G09_n, CGG, G09, RGG_n, G09_n, __A10_NET_204, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U10017(__A10_NET_206, __A10_NET_205, WHOMPA, __A10_2___XUY2, XUY10_n, __A10_NET_162, GND, __A10_1___RL_OUT_1, RLG_n, __A10_1___L1_n, GND, __A10_NET_202, G09, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U10018(__A10_NET_203, GND, SA09, __A10_NET_208, __A10_NET_207,  , GND,  , GND, SA10, __A10_NET_156, __A10_NET_155, __A10_NET_154, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10019(__A10_NET_150, A2XG_n, __A10_1___A2_n, __A10_NET_152, WYLOG_n, WL10_n, GND, WL09_n, WYDG_n, __A10_NET_151, __A10_1__Y2_n, CUG, __A10_1__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10020(MONEX, __A10_NET_150, __A10_1__X2_n, CLXC, CUG, __A10_1__X2, GND, __A10_1__Y2_n, __A10_NET_152, __A10_NET_151, __A10_1__Y2, __A10_1__X2_n, __A10_1__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10021(__A10_NET_144, __A10_1__X2_n, __A10_1__Y2_n, XUY10_n, __A10_1__X2, __A10_1__Y2, GND,  ,  ,  , __A10_NET_144, XUY10_n, __A10_NET_147, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10022( ,  , __A10_NET_144, __A10_1___SUMA2, CO10, __A10_2___CI_IN, GND, __A10_NET_148, __A10_1___SUMA2, __A10_1___SUMB2, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U10023(__A10_1___SUMB2, __A10_NET_147, __A10_NET_149, __A10_NET_133, WAG_n, WL10_n, GND, WL12_n, WALSG_n, __A10_NET_132, __A10_1___A2_n, CAG, __A10_NET_131, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10024(__A10_NET_133, __A10_NET_132, __A10_NET_148, __A10_NET_134, CH10, __A10_NET_129, GND, __A10_NET_139, __A10_NET_167, __A10_NET_168, __A10_NET_169, __A10_1___A2_n, __A10_NET_131, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10025(__A10_NET_134, RAG_n, __A10_1___A2_n, __A10_NET_167, WLG_n, WL10_n, GND, G13_n, G2LSG_n, __A10_NET_168, __A10_1___L2_n, CLG1G, __A10_NET_169, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10026(RLG_n, __A10_1___L2_n, __A10_1___RL_OUT_2, __A10_NET_135, __A10_NET_141, __A10_NET_140, GND, __A10_NET_130, MDT10, R1C, GND, __A10_1___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U10027(__A10_NET_171, WQG_n, WL10_n, __A10_1___Q2_n, __A10_NET_171, __A10_NET_170, GND, __A10_1___Q2_n, CQG, __A10_NET_170, RQG_n, __A10_1___Q2_n, __A10_NET_135, VCC, SIM_RST, SIM_CLK);
    assign RL10_n = RL10_n_U10028_2;
    assign __A10_1___Z2_n = __A10_1___Z2_n_U10028_4;
    assign RL10_n = RL10_n_U10028_6;
    assign RL10_n = RL10_n_U10028_8;
    assign G10_n = G10_n_U10028_10;
    assign G10_n = G10_n_U10028_12;
    U74LVC07 U10028(__A10_NET_140, RL10_n_U10028_2, __A10_NET_137, __A10_1___Z2_n_U10028_4, __A10_NET_130, RL10_n_U10028_6, GND, RL10_n_U10028_8, __A10_NET_172, G10_n_U10028_10, __A10_NET_154, G10_n_U10028_12, __A10_NET_161, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U10029(__A10_NET_136, WZG_n, WL10_n, __A10_NET_137, __A10_NET_136, __A10_NET_138, GND, __A10_1___Z2_n, CZG, __A10_NET_138, RZG_n, __A10_1___Z2_n, __A10_NET_141, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U10030(__A10_NET_175, WBG_n, WL10_n, __A10_1___B2_n, __A10_NET_175, __A10_NET_176, GND, __A10_1___B2_n, CBG, __A10_NET_176, RBLG_n, __A10_1___B2_n, __A10_NET_174, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U10031(__A10_NET_174, __A10_NET_173, __A10_NET_160, __A10_NET_159, G10, __A10_NET_161, GND, __A10_NET_255, GND, XUY14_n, __A10_2___XUY2, __A10_NET_172, __A10_NET_153, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10032(__A10_NET_173, __A10_NET_176, RCG_n, __A10_NET_156, WL09_n, WG3G_n, GND, WL11_n, WG4G_n, __A10_NET_155, L2GDG_n, __A10_1___L1_n, __A10_NET_160, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10033(__A10_NET_159, WG1G_n, WL10_n, G10, G10_n, CGG, GND, RGG_n, G10_n, __A10_NET_153,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U10034(G10_n, GEM10, RL10_n, __A10_1___WL2, __A10_1___WL2, WL10_n, GND, __A10_1___MWL2, RL10_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U10035(__A10_NET_290, A2XG_n, __A10_2___A1_n, __A10_NET_286, WYLOG_n, WL11_n, GND, WL10_n, WYDG_n, __A10_NET_285, __A10_2__Y1_n, CUG, __A10_2__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10036(MONEX, __A10_NET_290, __A10_2__X1_n, CLXC, CUG, __A10_2__X1, GND, __A10_2__Y1_n, __A10_NET_286, __A10_NET_285, __A10_2__Y1, __A10_2__X1_n, __A10_2__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10037(__A10_NET_294, __A10_2__X1_n, __A10_2__Y1_n, __A10_2___XUY1, __A10_2__X1, __A10_2__Y1, GND, __A10_NET_294, __A10_2___XUY1, __A10_NET_291, __A10_NET_294, SUMA11_n, __A10_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10038( ,  , SUMA11_n, SUMB11_n, RULOG_n, __A10_NET_272, GND, __A10_NET_276, XUY13_n, __A10_2___XUY1, __A10_2___CI_IN,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U10039(__A10_2___CI_IN, __A10_NET_292, G11_n, GEM11, RL11_n, __A10_2___WL1, GND, WL11_n, __A10_2___WL1, __A10_2___MWL1, RL11_n, __A10_NET_242, __A10_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10040(SUMB11_n, __A10_NET_291, __A10_NET_292, __A10_NET_275, WAG_n, WL11_n, GND, WL13_n, WALSG_n, __A10_NET_277, __A10_2___A1_n, CAG, __A10_NET_273, VCC, SIM_RST, SIM_CLK);
    assign CO14 = CO14_U10041_2;
    assign RL11_n = RL11_n_U10041_4;
    assign __A10_2___L1_n = __A10_2___L1_n_U10041_6;
    assign __A10_2___Z1_n = __A10_2___Z1_n_U10041_8;
    assign RL11_n = RL11_n_U10041_10;
    assign RL11_n = RL11_n_U10041_12;
    U74LVC07 U10041(__A10_NET_276, CO14_U10041_2, __A10_NET_271, RL11_n_U10041_4, __A10_NET_283, __A10_2___L1_n_U10041_6, GND, __A10_2___Z1_n_U10041_8, __A10_NET_306, RL11_n_U10041_10, __A10_NET_307, RL11_n_U10041_12, __A10_NET_305, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10042(__A10_NET_275, __A10_NET_277, __A10_NET_272, __A10_NET_270, CH11, __A10_NET_271, GND, __A10_NET_283, __A10_NET_274, __A10_NET_281, __A10_NET_282, __A10_2___A1_n, __A10_NET_273, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10043(__A10_NET_270, RAG_n, __A10_2___A1_n, __A10_NET_274, WLG_n, WL11_n, GND, G14_n, G2LSG_n, __A10_NET_281, __A10_2___L1_n, CLG1G, __A10_NET_282, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10044( ,  ,  ,  ,  ,  , GND, __A10_2___RL_OUT_1, RLG_n, __A10_2___L1_n, GND,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U10045( ,  ,  , __A10_NET_279, WQG_n, WL11_n, GND, __A10_NET_279, __A10_NET_278, __A10_2___Q1_n, __A10_2___Q1_n, CQG, __A10_NET_278, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U10046(__A10_NET_280, RQG_n, __A10_2___Q1_n, __A10_NET_309, WZG_n, WL11_n, GND, __A10_NET_309, __A10_NET_308, __A10_NET_306, __A10_2___Z1_n, CZG, __A10_NET_308, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U10047(__A10_NET_304, RZG_n, __A10_2___Z1_n, __A10_NET_313, WBG_n, WL11_n, GND, __A10_NET_313, __A10_NET_314, __A10_2___B1_n, __A10_2___B1_n, CBG, __A10_NET_314, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10048(__A10_NET_311, RBHG_n, __A10_2___B1_n, __A10_NET_312, __A10_NET_314, RCG_n, GND, WL10_n, WG3G_n, __A10_NET_301, WL12_n, WG4G_n, __A10_NET_300, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10049(__A10_2___RL_OUT_1, __A10_NET_280, MDT11, R1C, GND, __A10_NET_305, GND, __A10_NET_310, __A10_NET_311, __A10_NET_312, __A10_NET_297, __A10_NET_307, __A10_NET_304, VCC, SIM_RST, SIM_CLK);
    assign CO14 = CO14_U10050_2;
    assign RL11_n = RL11_n_U10050_4;
    assign G11_n = G11_n_U10050_6;
    assign G11_n = G11_n_U10050_8;
    assign RL12_n = RL12_n_U10050_10;
    assign L12_n = L12_n_U10050_12;
    U74LVC07 U10050(__A10_NET_255, CO14_U10050_2, __A10_NET_310, RL11_n_U10050_4, __A10_NET_296, G11_n_U10050_6, GND, G11_n_U10050_8, __A10_NET_295, RL12_n_U10050_10, __A10_NET_222, L12_n_U10050_12, __A10_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10051(__A10_NET_299, L2GDG_n, __A10_1___L2_n, __A10_NET_298, WG1G_n, WL11_n, GND, G11_n, CGG, G11, RGG_n, G11_n, __A10_NET_297, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U10052(__A10_NET_296, GND, SA11, __A10_NET_301, __A10_NET_300,  , GND,  , GND, SA12, __A10_NET_249, __A10_NET_248, __A10_NET_247, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U10053(__A10_NET_299, __A10_NET_298,  ,  ,  ,  , GND,  ,  ,  ,  , __A10_NET_295, G11, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10054(__A10_NET_243, A2XG_n, __A10_2___A2_n, __A10_NET_245, WYLOG_n, WL12_n, GND, WL11_n, WYDG_n, __A10_NET_244, __A10_2__Y2_n, CUG, __A10_2__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10055(MONEX, __A10_NET_243, __A10_2__X2_n, CLXC, CUG, __A10_2__X2, GND, __A10_2__Y2_n, __A10_NET_245, __A10_NET_244, __A10_2__Y2, __A10_2__X2_n, __A10_2__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10056(__A10_NET_237, __A10_2__X2_n, __A10_2__Y2_n, __A10_2___XUY2, __A10_2__X2, __A10_2__Y2, GND,  ,  ,  , __A10_NET_237, __A10_2___XUY2, __A10_NET_240, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10057( ,  , __A10_NET_237, SUMA12_n, __A10_2___CO_IN, CI13_n, GND, __A10_NET_241, SUMA12_n, SUMB12_n, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U10058(SUMB12_n, __A10_NET_240, __A10_NET_242, __A10_NET_226, WAG_n, WL12_n, GND, WL14_n, WALSG_n, __A10_NET_225, __A10_2___A2_n, CAG, __A10_NET_224, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10059(__A10_NET_226, __A10_NET_225, __A10_NET_241, __A10_NET_227, CH12, __A10_NET_222, GND, __A10_NET_232, __A10_NET_260, __A10_NET_261, __A10_NET_262, __A10_2___A2_n, __A10_NET_224, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10060(__A10_NET_227, RAG_n, __A10_2___A2_n, __A10_NET_260, WLG_n, WL12_n, GND, G15_n, G2LSG_n, __A10_NET_261, L12_n, CLG1G, __A10_NET_262, VCC, SIM_RST, SIM_CLK);
    U74HC27 U10061(RLG_n, L12_n, __A10_2___RL_OUT_2, __A10_NET_228, __A10_NET_234, __A10_NET_233, GND, __A10_NET_223, MDT12, R1C, GND, __A10_2___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U10062(__A10_NET_264, WQG_n, WL12_n, __A10_2___Q2_n, __A10_NET_264, __A10_NET_263, GND, __A10_2___Q2_n, CQG, __A10_NET_263, RQG_n, __A10_2___Q2_n, __A10_NET_228, VCC, SIM_RST, SIM_CLK);
    assign RL12_n = RL12_n_U10063_2;
    assign __A10_2___Z2_n = __A10_2___Z2_n_U10063_4;
    assign RL12_n = RL12_n_U10063_6;
    assign RL12_n = RL12_n_U10063_8;
    assign __A10_2___G2_n = __A10_2___G2_n_U10063_10;
    assign __A10_2___G2_n = __A10_2___G2_n_U10063_12;
    U74LVC07 U10063(__A10_NET_233, RL12_n_U10063_2, __A10_NET_230, __A10_2___Z2_n_U10063_4, __A10_NET_223, RL12_n_U10063_6, GND, RL12_n_U10063_8, __A10_NET_265, __A10_2___G2_n_U10063_10, __A10_NET_247, __A10_2___G2_n_U10063_12, __A10_NET_254, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U10064(__A10_NET_229, WZG_n, WL12_n, __A10_NET_230, __A10_NET_229, __A10_NET_231, GND, __A10_2___Z2_n, CZG, __A10_NET_231, RZG_n, __A10_2___Z2_n, __A10_NET_234, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U10065(__A10_NET_268, WBG_n, WL12_n, __A10_2___B2_n, __A10_NET_268, __A10_NET_269, GND, __A10_2___B2_n, CBG, __A10_NET_269, RBHG_n, __A10_2___B2_n, __A10_NET_267, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U10066(__A10_NET_267, __A10_NET_266, __A10_NET_253, __A10_NET_252, G12, __A10_NET_254, GND,  ,  ,  ,  , __A10_NET_265, __A10_NET_246, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10067(__A10_NET_266, __A10_NET_269, RCG_n, __A10_NET_249, WL11_n, WG3G_n, GND, WL13_n, WG4G_n, __A10_NET_248, L2GDG_n, __A10_2___L1_n, __A10_NET_253, VCC, SIM_RST, SIM_CLK);
    U74HC02 U10068(__A10_NET_252, WG1G_n, WL12_n, G12, __A10_2___G2_n, CGG, GND, RGG_n, __A10_2___G2_n, __A10_NET_246,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U10069(__A10_2___G2_n, GEM12, RL12_n, __A10_2___WL2, __A10_2___WL2, WL12_n, GND, __A10_2___MWL2, RL12_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC4002 U10070(__A10_1___SUMA1, __A10_NET_201, XUY09_n, CI09_n, GND,  , GND,  , __A10_NET_144, XUY10_n, __A10_1___CI_INTERNAL, GND, __A10_1___SUMA2, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U10071(SUMA11_n, __A10_NET_294, __A10_2___XUY1, __A10_2___CI_IN, GND,  , GND,  , __A10_NET_237, __A10_2___XUY2, __A10_2___CI_INTERNAL, WHOMP, SUMA12_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11001(__A11_NET_198, A2XG_n, __A11_1___A1_n, __A11_NET_193, WYHIG_n, WL13_n, GND, WL12_n, WYDG_n, __A11_NET_192, __A11_1__Y1_n, CUG, __A11_1__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11002(MONEX, __A11_NET_198, __A11_1__X1_n, CLXC, CUG, __A11_1__X1, GND, __A11_1__Y1_n, __A11_NET_193, __A11_NET_192, __A11_1__Y1, __A11_1__X1_n, __A11_1__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11003(__A11_NET_202, __A11_1__X1_n, __A11_1__Y1_n, XUY13_n, __A11_1__X1, __A11_1__Y1, GND, __A11_NET_202, XUY13_n, __A11_NET_200, __A11_NET_202, SUMA13_n, __A11_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11004( ,  , SUMA13_n, SUMB13_n, RULOG_n, __A11_NET_180, GND, __A11_NET_184, __A11_2___XUY1, XUY13_n, CI13_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U11005(CI13_n, __A11_NET_199, G13_n, GEM13, RL13_n, __A11_1___WL1, GND, WL13_n, __A11_1___WL1, __A11_1___MWL1, RL13_n, __A11_NET_150, __A11_1___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11006(SUMB13_n, __A11_NET_200, __A11_NET_199, __A11_NET_183, WAG_n, WL13_n, GND, WL15_n, WALSG_n, __A11_NET_185, __A11_1___A1_n, CAG, __A11_NET_181, VCC, SIM_RST, SIM_CLK);
    assign __A11_2___CO_IN = __A11_2___CO_IN_U11007_2;
    assign RL13_n = RL13_n_U11007_4;
    assign __A11_1___L1_n = __A11_1___L1_n_U11007_6;
    assign __A11_1___Z1_n = __A11_1___Z1_n_U11007_8;
    assign RL13_n = RL13_n_U11007_10;
    assign RL13_n = RL13_n_U11007_12;
    U74LVC07 U11007(__A11_NET_184, __A11_2___CO_IN_U11007_2, __A11_NET_178, RL13_n_U11007_4, __A11_NET_191, __A11_1___L1_n_U11007_6, GND, __A11_1___Z1_n_U11007_8, __A11_NET_214, RL13_n_U11007_10, __A11_NET_215, RL13_n_U11007_12, __A11_NET_213, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11008(__A11_NET_179, RAG_n, __A11_1___A1_n, __A11_NET_182, WLG_n, WL13_n, GND, WL01_n, WALSG_n, __A11_NET_189, __A11_1___L1_n, CLG2G, __A11_NET_190, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11009( ,  ,  , __A11_NET_187, WQG_n, WL13_n, GND, __A11_NET_187, __A11_NET_186, __A11_1___Q1_n, __A11_1___Q1_n, CQG, __A11_NET_186, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11010(__A11_NET_188, RQG_n, __A11_1___Q1_n, __A11_NET_217, WZG_n, WL13_n, GND, __A11_NET_217, __A11_NET_216, __A11_NET_214, __A11_1___Z1_n, CZG, __A11_NET_216, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11011(__A11_1___RL_OUT_1, __A11_NET_188, MDT13, R1C, GND, __A11_NET_213, GND, __A11_NET_220, __A11_NET_218, __A11_NET_219, __A11_NET_205, __A11_NET_215, __A11_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11012(__A11_NET_212, RZG_n, __A11_1___Z1_n, __A11_NET_221, WBG_n, WL13_n, GND, __A11_NET_221, __A11_NET_222, __A11_1___B1_n, __A11_1___B1_n, CBG, __A11_NET_222, VCC, SIM_RST, SIM_CLK);
    assign __A11_2___CO_IN = __A11_2___CO_IN_U11013_2;
    assign RL13_n = RL13_n_U11013_4;
    assign G13_n = G13_n_U11013_6;
    assign G13_n = G13_n_U11013_8;
    assign RL14_n = RL14_n_U11013_10;
    assign __A11_1___L2_n = __A11_1___L2_n_U11013_12;
    U74LVC07 U11013(__A11_NET_163, __A11_2___CO_IN_U11013_2, __A11_NET_220, RL13_n_U11013_4, __A11_NET_204, G13_n_U11013_6, GND, G13_n_U11013_8, __A11_NET_203, RL14_n_U11013_10, __A11_NET_130, __A11_1___L2_n_U11013_12, __A11_NET_140, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11014(__A11_NET_218, RBHG_n, __A11_1___B1_n, __A11_NET_219, __A11_NET_222, RCG_n, GND, WL12_n, WG3G_n, __A11_NET_209, WL14_n, WG4G_n, __A11_NET_208, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11015(__A11_NET_183, __A11_NET_185, __A11_NET_180, __A11_NET_179, CH13, __A11_NET_178, GND, __A11_NET_191, __A11_NET_182, __A11_NET_189, __A11_NET_190, __A11_1___A1_n, __A11_NET_181, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11016(__A11_NET_207, L2GDG_n, L12_n, __A11_NET_206, WG1G_n, WL13_n, GND, G13_n, CGG, G13, RGG_n, G13_n, __A11_NET_205, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U11017(__A11_NET_207, __A11_NET_206, GND, __A11_2___XUY2, XUY14_n, __A11_NET_163, GND, __A11_1___RL_OUT_1, RLG_n, __A11_1___L1_n, GND, __A11_NET_203, G13, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U11018(__A11_NET_204, GND, SA13, __A11_NET_209, __A11_NET_208,  , GND,  , GND, SA14, __A11_NET_157, __A11_NET_156, __A11_NET_155, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11019(__A11_NET_151, A2XG_n, __A11_1___A2_n, __A11_NET_153, WYHIG_n, WL14_n, GND, WL13_n, WYDG_n, __A11_NET_152, __A11_1__Y2_n, CUG, __A11_1__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11020(MONEX, __A11_NET_151, __A11_1__X2_n, CLXC, CUG, __A11_1__X2, GND, __A11_1__Y2_n, __A11_NET_153, __A11_NET_152, __A11_1__Y2, __A11_1__X2_n, __A11_1__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11021(__A11_NET_145, __A11_1__X2_n, __A11_1__Y2_n, XUY14_n, __A11_1__X2, __A11_1__Y2, GND,  ,  ,  , __A11_NET_145, XUY14_n, __A11_NET_148, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11022( ,  , __A11_NET_145, SUMA14_n, CO14, __A11_2___CI_IN, GND, __A11_NET_149, SUMA14_n, SUMB14_n, RULOG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U11023(SUMB14_n, __A11_NET_148, __A11_NET_150, __A11_NET_134, WAG_n, WL14_n, GND, WL16_n, WALSG_n, __A11_NET_133, __A11_1___A2_n, CAG, __A11_NET_132, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11024(__A11_NET_134, __A11_NET_133, __A11_NET_149, __A11_NET_135, CH14, __A11_NET_130, GND, __A11_NET_140, __A11_NET_168, __A11_NET_169, __A11_NET_170, __A11_1___A2_n, __A11_NET_132, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11025(__A11_NET_135, RAG_n, __A11_1___A2_n, __A11_NET_168, WLG_n, WL14_n, GND, WL02_n, WALSG_n, __A11_NET_169, __A11_1___L2_n, CLG2G, __A11_NET_170, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11026(RLG_n, __A11_1___L2_n, __A11_1___RL_OUT_2, __A11_NET_136, __A11_NET_142, __A11_NET_141, GND, __A11_NET_131, MDT14, R1C, GND, __A11_1___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11027(__A11_NET_172, WQG_n, WL14_n, __A11_1___Q2_n, __A11_NET_172, __A11_NET_171, GND, __A11_1___Q2_n, CQG, __A11_NET_171, RQG_n, __A11_1___Q2_n, __A11_NET_136, VCC, SIM_RST, SIM_CLK);
    assign RL14_n = RL14_n_U11028_2;
    assign __A11_1___Z2_n = __A11_1___Z2_n_U11028_4;
    assign RL14_n = RL14_n_U11028_6;
    assign RL14_n = RL14_n_U11028_8;
    assign G14_n = G14_n_U11028_10;
    assign G14_n = G14_n_U11028_12;
    U74LVC07 U11028(__A11_NET_141, RL14_n_U11028_2, __A11_NET_138, __A11_1___Z2_n_U11028_4, __A11_NET_131, RL14_n_U11028_6, GND, RL14_n_U11028_8, __A11_NET_173, G14_n_U11028_10, __A11_NET_155, G14_n_U11028_12, __A11_NET_162, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11029(__A11_NET_137, WZG_n, WL14_n, __A11_NET_138, __A11_NET_137, __A11_NET_139, GND, __A11_1___Z2_n, CZG, __A11_NET_139, RZG_n, __A11_1___Z2_n, __A11_NET_142, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11030(__A11_NET_176, WBG_n, WL14_n, __A11_1___B2_n, __A11_NET_176, __A11_NET_177, GND, __A11_1___B2_n, CBG, __A11_NET_177, RBHG_n, __A11_1___B2_n, __A11_NET_175, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U11031(__A11_NET_175, __A11_NET_174, __A11_NET_161, __A11_NET_160, G14, __A11_NET_162, GND, __A11_NET_256, GND, XUY02_n, __A11_2___XUY2, __A11_NET_173, __A11_NET_154, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11032(__A11_NET_174, __A11_NET_177, RCG_n, __A11_NET_157, WL13_n, WG3G_n, GND, WL16_n, WG4G_n, __A11_NET_156, L2GDG_n, __A11_1___L1_n, __A11_NET_161, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11033(__A11_NET_160, WG1G_n, WL14_n, G14, G14_n, CGG, GND, RGG_n, G14_n, __A11_NET_154,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U11034(G14_n, GEM14, RL14_n, __A11_1___WL2, __A11_1___WL2, WL14_n, GND, __A11_1___MWL2, RL14_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U11035(__A11_NET_291, A2XG_n, __A11_2___A1_n, __A11_NET_287, WYHIG_n, WL15_n, GND, WL14_n, WYDG_n, __A11_NET_286, __A11_2__Y1_n, CUG, __A11_2__Y1, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11036(BXVX, __A11_NET_291, __A11_2__X1_n, CLXC, CUG, __A11_2__X1, GND, __A11_2__Y1_n, __A11_NET_287, __A11_NET_286, __A11_2__Y1, __A11_2__X1_n, __A11_2__X1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11037(__A11_NET_295, __A11_2__X1_n, __A11_2__Y1_n, __A11_2___XUY1, __A11_2__X1, __A11_2__Y1, GND, __A11_NET_295, __A11_2___XUY1, __A11_NET_292, __A11_NET_295, SUMA15_n, __A11_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11038( ,  , SUMA15_n, SUMB15_n, RULOG_n, __A11_NET_273, GND, __A11_NET_277, XUY01_n, __A11_2___XUY1, __A11_2___CI_IN,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U11039(__A11_2___CI_IN, __A11_NET_293, G15_n, __A11_2___GEM1, RL15_n, WL15, GND, WL15_n, WL15, __A11_2___MWL1, RL15_n, __A11_NET_243, __A11_2___CI_INTERNAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11040(SUMB15_n, __A11_NET_292, __A11_NET_293, __A11_NET_276, WAG_n, WL15_n, GND, G16SW_n, WALSG_n, __A11_NET_278, __A11_2___A1_n, CAG, __A11_NET_274, VCC, SIM_RST, SIM_CLK);
    assign __A11_2___CO_OUT = __A11_2___CO_OUT_U11041_2;
    assign RL15_n = RL15_n_U11041_4;
    assign L15_n = L15_n_U11041_6;
    assign Z15_n = Z15_n_U11041_8;
    assign RL15_n = RL15_n_U11041_10;
    assign RL15_n = RL15_n_U11041_12;
    U74LVC07 U11041(__A11_NET_277, __A11_2___CO_OUT_U11041_2, __A11_NET_272, RL15_n_U11041_4, __A11_NET_284, L15_n_U11041_6, GND, Z15_n_U11041_8, __A11_NET_307, RL15_n_U11041_10, __A11_NET_308, RL15_n_U11041_12, __A11_NET_306, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11042(__A11_NET_276, __A11_NET_278, __A11_NET_273, __A11_NET_271, CH16, __A11_NET_272, GND, __A11_NET_284, __A11_NET_275, __A11_NET_282, __A11_NET_283, __A11_2___A1_n, __A11_NET_274, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11043(__A11_NET_271, RAG_n, __A11_2___A1_n, __A11_NET_275, WLG_n, WL15_n, GND, G01_n, G2LSG_n, __A11_NET_282, L15_n, CLG1G, __A11_NET_283, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11044( ,  ,  ,  ,  ,  , GND, __A11_2___RL_OUT_1, RLG_n, L15_n, VCC,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11045( ,  ,  , __A11_NET_280, WQG_n, WL15_n, GND, __A11_NET_280, __A11_NET_279, __A11_2___Q1_n, __A11_2___Q1_n, CQG, __A11_NET_279, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11046(__A11_NET_281, RQG_n, __A11_2___Q1_n, __A11_NET_310, WZG_n, WL15_n, GND, __A11_NET_310, __A11_NET_309, __A11_NET_307, Z15_n, CZG, __A11_NET_309, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11047(__A11_NET_305, RZG_n, Z15_n, __A11_NET_314, WBG_n, WL15_n, GND, __A11_NET_314, __A11_NET_315, __A11_2___B1_n, __A11_2___B1_n, CBG, __A11_NET_315, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11048(__A11_NET_312, RBHG_n, __A11_2___B1_n, __A11_NET_313, __A11_NET_315, RCG_n, GND, GND, VCC, __A11_NET_302, GND, VCC, __A11_NET_301, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11049(__A11_2___RL_OUT_1, __A11_NET_281, MDT15, R1C, __A11_2___RL_OUT_2, __A11_NET_306, GND, __A11_NET_311, __A11_NET_312, __A11_NET_313, __A11_NET_298, __A11_NET_308, __A11_NET_305, VCC, SIM_RST, SIM_CLK);
    assign __A11_2___CO_OUT = __A11_2___CO_OUT_U11050_2;
    assign RL15_n = RL15_n_U11050_4;
    assign G15_n = G15_n_U11050_6;
    assign G15_n = G15_n_U11050_8;
    assign RL16_n = RL16_n_U11050_10;
    assign L16_n = L16_n_U11050_12;
    U74LVC07 U11050(__A11_NET_256, __A11_2___CO_OUT_U11050_2, __A11_NET_311, RL15_n_U11050_4, __A11_NET_297, G15_n_U11050_6, GND, G15_n_U11050_8, __A11_NET_296, RL16_n_U11050_10, __A11_NET_223, L16_n_U11050_12, __A11_NET_233, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11051(__A11_NET_300, L2GDG_n, __A11_1___L2_n, __A11_NET_299, WG1G_n, WL15_n, GND, G15_n, CGG, G15, RGG_n, G15_n, __A11_NET_298, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U11052(__A11_NET_297, GND, SA16, __A11_NET_302, __A11_NET_301,  , GND,  , GND, SA16, __A11_NET_250, __A11_NET_249, __A11_NET_248, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U11053(__A11_NET_300, __A11_NET_299,  ,  ,  ,  , GND,  ,  ,  ,  , __A11_NET_296, G15, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11054(__A11_NET_244, A2XG_n, __A11_2___A2_n, __A11_NET_246, WYHIG_n, WL16_n, GND, WL16_n, WYDG_n, __A11_NET_245, __A11_2__Y2_n, CUG, __A11_2__Y2, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11055(MONEX, __A11_NET_244, __A11_2__X2_n, CLXC, CUG, __A11_2__X2, GND, __A11_2__Y2_n, __A11_NET_246, __A11_NET_245, __A11_2__Y2, __A11_2__X2_n, __A11_2__X2, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11056(__A11_NET_238, __A11_2__X2_n, __A11_2__Y2_n, __A11_2___XUY2, __A11_2__X2, __A11_2__Y2, GND,  ,  ,  , __A11_NET_238, __A11_2___XUY2, __A11_NET_241, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11057( ,  , __A11_NET_238, SUMA16_n, __A11_2___CO_IN, EAC_n, GND, __A11_NET_242, SUMA16_n, SUMB16_n, RUG_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U11058(SUMB16_n, __A11_NET_241, __A11_NET_243, __A11_NET_227, WAG_n, WL16_n, GND, G16SW_n, WALSG_n, __A11_NET_226, __A11_2___A2_n, CAG, __A11_NET_225, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11059(__A11_NET_227, __A11_NET_226, __A11_NET_242, __A11_NET_228, CH16, __A11_NET_223, GND, __A11_NET_233, __A11_NET_261, __A11_NET_262, __A11_NET_263, __A11_2___A2_n, __A11_NET_225, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11060(__A11_NET_228, RAG_n, __A11_2___A2_n, __A11_NET_261, WLG_n, WL16_n, GND, __A11_2___G2_n, G2LSG_n, __A11_NET_262, L16_n, CLG1G, __A11_NET_263, VCC, SIM_RST, SIM_CLK);
    U74HC27 U11061(RLG_n, L16_n, __A11_2___RL_OUT_2, __A11_NET_229, __A11_NET_235, __A11_NET_234, GND, __A11_NET_224, MDT16, R1C, US2SG, __A11_2___RL_OUT_2, GND, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11062(__A11_NET_265, WQG_n, WL16_n, __A11_2___Q2_n, __A11_NET_265, __A11_NET_264, GND, __A11_2___Q2_n, CQG, __A11_NET_264, RQG_n, __A11_2___Q2_n, __A11_NET_229, VCC, SIM_RST, SIM_CLK);
    assign RL16_n = RL16_n_U11063_2;
    assign Z16_n = Z16_n_U11063_4;
    assign RL16_n = RL16_n_U11063_6;
    assign RL16_n = RL16_n_U11063_8;
    assign __A11_2___G2_n = __A11_2___G2_n_U11063_10;
    assign __A11_2___G2_n = __A11_2___G2_n_U11063_12;
    U74LVC07 U11063(__A11_NET_234, RL16_n_U11063_2, __A11_NET_231, Z16_n_U11063_4, __A11_NET_224, RL16_n_U11063_6, GND, RL16_n_U11063_8, __A11_NET_266, __A11_2___G2_n_U11063_10, __A11_NET_248, __A11_2___G2_n_U11063_12, __A11_NET_255, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11064(__A11_NET_230, WZG_n, WL16_n, __A11_NET_231, __A11_NET_230, __A11_NET_232, GND, Z16_n, CZG, __A11_NET_232, RZG_n, Z16_n, __A11_NET_235, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11065(__A11_NET_269, WBG_n, WL16_n, __A11_2___B2_n, __A11_NET_269, __A11_NET_270, GND, __A11_2___B2_n, CBG, __A11_NET_270, RBHG_n, __A11_2___B2_n, __A11_NET_268, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U11066(__A11_NET_268, __A11_NET_267, __A11_NET_254, __A11_NET_253, G16, __A11_NET_255, GND,  ,  ,  ,  , __A11_NET_266, __A11_NET_247, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11067(__A11_NET_267, __A11_NET_270, RCG_n, __A11_NET_250, WL14_n, WG3G_n, GND, WL01_n, WG5G_n, __A11_NET_249, L2GDG_n, L16_n, __A11_NET_254, VCC, SIM_RST, SIM_CLK);
    U74HC02 U11068(__A11_NET_253, WG2G_n, WL16_n, G16, __A11_2___G2_n, CGG, GND, RGG_n, __A11_2___G2_n, __A11_NET_247,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U11069(__A11_2___G2_n, GEM16, RL16_n, WL16, WL16, WL16_n, GND, __A11_2___MWL2, RL16_n,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC4002 U11070(SUMA13_n, __A11_NET_202, XUY13_n, CI13_n, GND,  , GND,  , __A11_NET_145, XUY14_n, __A11_1___CI_INTERNAL, GND, SUMA14_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U11071(SUMA15_n, __A11_NET_295, __A11_2___XUY1, __A11_2___CI_IN, GND,  , GND,  , __A11_NET_238, __A11_2___XUY2, __A11_2___CI_INTERNAL, WHOMPA, SUMA16_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12001(G01, __A12_1__G01A_n, G02, __A12_1__G02_n, G03, __A12_1__G03_n, GND, __A12_1__PA03_n, __A12_1__PA03, __A12_NET_198, G04, __A12_NET_191, G05, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12002(G01, G02, G01, __A12_1__G02_n, __A12_1__G03_n, __A12_NET_181, GND, __A12_NET_185, __A12_1__G01A_n, G02, __A12_1__G03_n, __A12_NET_180, G03, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12003(__A12_1__G01A_n, __A12_1__G02_n, G04, G05, G06, __A12_NET_186, GND, __A12_NET_192, G04, __A12_NET_191, __A12_NET_197, __A12_NET_184, G03, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U12004(__A12_1__PA03, __A12_NET_180, __A12_NET_181, __A12_NET_185, __A12_NET_184,  , GND,  , __A12_NET_186, __A12_NET_192, __A12_NET_190, __A12_NET_187, __A12_1__PA06, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12005(G06, __A12_NET_197, __A12_NET_186, __A12_NET_139, __A12_1__PA06, __A12_1__PA06_n, GND, __A12_NET_196, G07, __A12_NET_131, G08, __A12_NET_177, G09, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12006(__A12_NET_198, G05, __A12_NET_198, __A12_NET_191, G06, __A12_NET_187, GND, __A12_NET_127, G07, G08, G09, __A12_NET_190, __A12_NET_197, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12007(G07, __A12_NET_131, __A12_NET_196, G08, __A12_NET_177, __A12_NET_129, GND, __A12_NET_128, __A12_NET_196, __A12_NET_131, G09, __A12_NET_125, __A12_NET_177, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U12008(__A12_1__PA09, __A12_NET_127, __A12_NET_125, __A12_NET_129, __A12_NET_128,  , GND,  , __A12_NET_141, __A12_NET_130, __A12_NET_143, __A12_NET_142, __A12_1__PA12, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12009(__A12_NET_127, __A12_NET_138, __A12_1__PA09, __A12_1__PA09_n, G10, __A12_NET_124, GND, __A12_NET_126, G11, __A12_NET_123, G12, __A12_NET_137, __A12_NET_141, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12010(G10, G11, G10, __A12_NET_126, __A12_NET_123, __A12_NET_130, GND, __A12_NET_143, __A12_NET_124, G11, __A12_NET_123, __A12_NET_141, G12, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12011(__A12_NET_124, __A12_NET_126, G13, G14, G16, __A12_NET_135, GND, __A12_NET_134, G13, __A12_NET_136, __A12_1__G16A_n, __A12_NET_142, G12, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12012(__A12_1__PA12, __A12_1__PA12_n, G13, __A12_NET_140, G14, __A12_NET_136, GND, __A12_1__G16A_n, G16, __A12_NET_117, __A12_NET_135, __A12_1__PA15_n, __A12_1__PA15, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12013(__A12_NET_140, G14, __A12_NET_140, __A12_NET_136, G16, __A12_NET_132, GND, __A12_NET_199, __A12_NET_139, __A12_NET_138, __A12_NET_137, __A12_NET_133, __A12_1__G16A_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b0, 1'b1) U12014(__A12_1__PA15, __A12_NET_135, __A12_NET_134, __A12_NET_133, __A12_NET_132,  , GND,  , EXTPLS, RELPLS, INHPLS, __A12_NET_122, __A12_NET_121, VCC, SIM_RST, SIM_CLK);
    U74HC02 U12015(__A12_NET_200, __A12_NET_117, G15, __A12_NET_114, TSUDO_n, __A12_1__T7PHS4_n, GND, __A12_1__G02_n, G03, __A12_NET_195, G02, __A12_1__G03_n, __A12_NET_193, VCC, SIM_RST, SIM_CLK);
    assign __A12_1__GNZRO = __A12_1__GNZRO_U12016_2;
    assign __A12_1__GNZRO = __A12_1__GNZRO_U12016_4;
    assign RELPLS = RELPLS_U12016_6;
    assign RELPLS = RELPLS_U12016_8;
    assign INHPLS = INHPLS_U12016_10;
    assign INHPLS = INHPLS_U12016_12;
    U74LVC07 U12016(__A12_NET_199, __A12_1__GNZRO_U12016_2, __A12_NET_200, __A12_1__GNZRO_U12016_4, __A12_NET_201, RELPLS_U12016_6, GND, RELPLS_U12016_8, __A12_NET_195, INHPLS_U12016_10, __A12_NET_194, INHPLS_U12016_12, __A12_NET_193, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12017(__A12_1__GNZRO, __A12_NET_115, __A12_NET_181, __A12_NET_116, __A12_NET_114, __A12_NET_113, GND, GEQZRO_n, __A12_NET_110, __A12_NET_119, RAD, __A12_1__PB09_n, __A12_1__PB09, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12018(__A12_NET_116, __A12_NET_115, __A12_NET_115, __A12_NET_113, __A12_1__G01A_n, __A12_NET_201, GND, __A12_NET_194, __A12_NET_115, G01, __A12_NET_113, EXTPLS, __A12_NET_113, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U12019(__A12_NET_110, __A12_NET_115, G02, G01, G03,  , GND,  , __A12_NET_155, __A12_NET_154, __A12_NET_153, __A12_NET_163, __A12_1__PB09, VCC, SIM_RST, SIM_CLK);
    U74HC02 U12020(__A12_NET_122, __A12_NET_121, T12A, RADRZ, __A12_NET_121, __A12_NET_119, GND, __A12_NET_119, __A12_NET_122, RADRG, __A12_1__PA12, __A12_1__PA15, __A12_NET_152, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12021(__A12_1__PA03, __A12_1__PA06, __A12_1__PA03, __A12_1__PA06_n, __A12_1__PA09_n, __A12_NET_154, GND, __A12_NET_153, __A12_1__PA03_n, __A12_1__PA06, __A12_1__PA09_n, __A12_NET_155, __A12_1__PA09, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U12022(__A12_1__PA03_n, __A12_1__PA06_n, __A12_NET_145, MONPAR, SAP, __A12_NET_146, GND, __A12_NET_144, SCAD, __A12_NET_147, GOJAM, __A12_NET_163, __A12_1__PA09, VCC, SIM_RST, SIM_CLK);
    U74HC02 U12023(__A12_NET_158, __A12_1__PA12_n, __A12_1__PA15_n, __A12_1__PB15, __A12_NET_152, __A12_NET_158, GND, __A12_1__PB09_n, __A12_1__PB15, __A12_NET_170, __A12_1__PB09, __A12_1__PB15_n, __A12_NET_171, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12024(__A12_1__PB15, __A12_1__PB15_n, __A12_1__PC15, PC15_n, __A12_1__PC15, __A12_1__MGP_n, GND, GEMP, PC15_n, __A12_1__MSP, __A12_NET_146, __A12_1__MPAL, PALE, VCC, SIM_RST, SIM_CLK);
    U74HC02 U12025(__A12_1__PC15, __A12_NET_170, __A12_NET_171, __A12_NET_145, CGG, __A12_NET_146, GND, __A12_1__PC15, __A12_NET_145, __A12_NET_147, PC15_n, __A12_NET_146, __A12_NET_150, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12026(TPARG_n, n8XP5, T07_n, PHS4_n, FUTEXT, __A12_1__T7PHS4, GND, __A12_NET_243, XB0_n, T02_n, __A12_NET_245, __A12_NET_151, __A12_NET_150, VCC, SIM_RST, SIM_CLK);
    assign PALE = PALE_U12027_2;
    assign PALE = PALE_U12027_4;
    U74LVC07 U12027(__A12_NET_144, PALE_U12027_2, __A12_NET_151, PALE_U12027_4,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12028(G01ED, WEDOPG_n, WL08_n, __A12_NET_256, WL08_n, WSG_n, GND, __A12_NET_256, __A12_NET_235, __A12_NET_257, __A12_NET_257, CSG, __A12_NET_235, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12029(__A12_NET_257, S08, __A12_NET_235, S08_n, __A12_NET_237, S09, GND, S09_n, __A12_NET_236, S10, __A12_NET_229, S10_n, __A12_NET_230, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12030(G02ED, WEDOPG_n, WL09_n, __A12_NET_238, WL09_n, WSG_n, GND, __A12_NET_238, __A12_NET_236, __A12_NET_237, __A12_NET_237, CSG, __A12_NET_236, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12031(G03ED, WEDOPG_n, WL10_n, __A12_NET_239, WL10_n, WSG_n, GND, __A12_NET_239, __A12_NET_230, __A12_NET_229, __A12_NET_229, CSG, __A12_NET_230, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12032(G04ED, WEDOPG_n, WL11_n, __A12_NET_228, WL11_n, WSG_n, GND, __A12_NET_228, __A12_NET_231, __A12_NET_232, __A12_NET_232, CSG, __A12_NET_231, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12033(__A12_NET_232, S11, __A12_NET_231, S11_n, __A12_NET_234, S12, GND, S12_n, __A12_NET_233, S01, __A12_NET_227, S01_n, __A12_NET_226, VCC, SIM_RST, SIM_CLK);
    U74HC02 U12034(G05ED, WEDOPG_n, WL12_n, __A12_NET_241, WL12_n, WSG_n, GND, EDOP_n, T12A, __A12_NET_251, __A12_NET_234, CSG, __A12_NET_233, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U12035(G06ED, WEDOPG_n, WL13_n, G07ED, WEDOPG_n, WL14_n, GND, WL01_n, WSG_n, __A12_NET_240, __A12_NET_240, __A12_NET_226, __A12_NET_227, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12036(__A12_NET_226, __A12_NET_227, CSG, __A12_NET_217, WL02_n, WSG_n, GND, __A12_NET_217, __A12_NET_218, __A12_NET_219, __A12_NET_219, CSG, __A12_NET_218, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12037(__A12_NET_219, S02, __A12_NET_218, S02_n, __A12_NET_221, S03, GND, S03_n, __A12_NET_216, S04, __A12_NET_211, S04_n, __A12_NET_210, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U12038(__A12_NET_220, WL03_n, WSG_n, __A12_NET_221, __A12_NET_220, __A12_NET_216, GND, __A12_NET_221, CSG, __A12_NET_216, WL04_n, WSG_n, __A12_NET_222, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U12039(__A12_NET_211, __A12_NET_222, __A12_NET_210, __A12_NET_210, __A12_NET_211, CSG, GND, WL05_n, WSG_n, __A12_NET_209, __A12_NET_209, __A12_NET_208, __A12_NET_207, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12040(__A12_NET_208, __A12_NET_207, CSG, __A12_NET_212, WL06_n, WSG_n, GND, __A12_NET_212, __A12_NET_213, __A12_NET_214, __A12_NET_214, CSG, __A12_NET_213, VCC, SIM_RST, SIM_CLK);
    U74HC04 U12041(__A12_NET_207, S05, __A12_NET_208, S05_n, __A12_NET_214, S06, GND, S06_n, __A12_NET_213, S07, __A12_NET_224, S07_n, __A12_NET_225, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U12042(__A12_NET_215, WL07_n, WSG_n, __A12_NET_224, __A12_NET_215, __A12_NET_225, GND, __A12_NET_224, CSG, __A12_NET_225,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U12043(__A12_1__T7PHS4, __A12_1__T7PHS4_n,  ,  , OCTAD2, __A12_NET_245, GND, GINH, __A12_NET_223, __A12_2__G01A, __A12_1__G01A_n,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC4002 U12044( ,  ,  ,  ,  ,  , GND,  , __A12_NET_242, __A12_NET_244, __A12_NET_254, __A12_NET_251, __A12_NET_223, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U12046( ,  ,  , CYR_n, __A12_NET_243, __A12_NET_242, GND, CYR_n, T12A, __A12_NET_242, __A12_NET_246, __A12_NET_244, SR_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U12047(__A12_NET_245, T02_n, __A12_NET_245, T02_n, XB2_n, __A12_NET_255, GND, __A12_NET_250, __A12_NET_245, T02_n, XB3_n, __A12_NET_246, XB1_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U12048(__A12_NET_244, SR_n, T12A, CYL_n, __A12_NET_255, __A12_NET_254, GND, CYL_n, T12A, __A12_NET_254, __A12_NET_250, __A12_NET_251, EDOP_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U12049(n8XP5, __A12_NET_241, SUMA16_n, SUMB16_n, __A12_1__G01A_n, __A12_NET_248, GND,  ,  ,  ,  , __A12_NET_234, __A12_NET_233, VCC, SIM_RST, SIM_CLK);
    U74HC02 U12050(__A12_NET_249, __A12_2__G01A, __A12_1__G16A_n, G16SW_n, __A12_NET_249, __A12_NET_248, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U13001(MSTRT, __A13_NET_235, F12B, __A13_1__F12B_n, __A13_1__F14H, __A13_NET_221, GND, __A13_NET_265, __A13_NET_266, __A13_1__NOTEST, __A13_1__NOTEST_n, __A13_1__DOFILT, __A13_NET_254, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U13002(__A13_NET_238, F05B_n, __A13_NET_235, __A13_NET_236, __A13_NET_238, __A13_NET_237, GND, __A13_NET_236, __A13_NET_235, __A13_NET_237, F05A_n, __A13_NET_236, MSTRTP, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U13003(__A13_NET_233, IIP, __A13_NET_222, __A13_NET_222, __A13_NET_233, F14B, GND, IIP_n, __A13_NET_223, __A13_NET_226, __A13_NET_226, F14B, __A13_NET_223, VCC, SIM_RST, SIM_CLK);
    U74HC27 U13004(__A13_1__F12B_n, FS14, PALE, __A13_NET_230, __A13_NET_229, __A13_NET_249, GND, __A13_NET_250, __A13_NET_244, __A13_NET_231, __A13_1__WATCHP, __A13_1__F14H, __A13_1__FS13_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U13005(__A13_NET_230, __A13_NET_222, __A13_NET_221, __A13_NET_229, __A13_NET_223, __A13_NET_221, GND, __A13_NET_230, __A13_NET_229, __A13_1__MRPTAL_n, __A13_NET_228, F10B, __A13_NET_232, VCC, SIM_RST, SIM_CLK);
    assign __A13_1__CKTAL_n = __A13_1__CKTAL_n_U13006_2;
    assign __A13_1__CKTAL_n = __A13_1__CKTAL_n_U13006_4;
    assign __A13_NET_266 = __A13_NET_266_U13006_6;
    assign __A13_NET_266 = __A13_NET_266_U13006_8;
    assign __A13_NET_266 = __A13_NET_266_U13006_10;
    assign __A13_NET_266 = __A13_NET_266_U13006_12;
    U74LVC07 U13006(__A13_NET_249, __A13_1__CKTAL_n_U13006_2, __A13_NET_250, __A13_1__CKTAL_n_U13006_4, __A13_NET_206, __A13_NET_266_U13006_6, GND, __A13_NET_266_U13006_8, __A13_NET_192, __A13_NET_266_U13006_10, __A13_NET_193, __A13_NET_266_U13006_12, __A13_NET_187, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U13007(TC0, TCF0, T12_n, PHS4_n, NISQL_n, __A13_NET_298, GND, __A13_NET_270, __A13_1__NOTEST, __A13_NET_263, T09_n, __A13_NET_228, __A13_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U13008(__A13_NET_234, __A13_NET_243, __A13_NET_227, __A13_NET_227, __A13_NET_234, F10B, GND, __A13_NET_232, F10A_n, __A13_NET_244, __A13_NET_227, F10A_n, __A13_NET_231, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U13009(__A13_NET_243, TCF0, TC0, INKL, T04_n,  , GND,  , INLNKP, INLNKM, RNRADP, RNRADM, __A13_NET_199, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U13010(__A13_1__MTCAL_n, __A13_NET_244, __A13_NET_231, __A13_NET_263, __A13_NET_265, __A13_NET_264, GND, __A13_NET_263, INKL, __A13_NET_264, PSEUDO, NISQL_n, __A13_1__NOTEST_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U13011(__A13_NET_198, GYROD, CDUXD, CDUYD, CDUZD,  , GND,  , TRUND, SHAFTD, THRSTD, EMSD, __A13_NET_197, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U13012(__A13_NET_273, __A13_NET_270, __A13_NET_272, __A13_NET_272, __A13_NET_273, INKL, GND, T03_n, __A13_NET_273, __A13_NET_253, __A13_NET_253, __A13_NET_257, __A13_1__MCTRAL_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U13013(INKL, T03_n, __A13_NET_253, __A13_NET_257, GOJAM, __A13_NET_254, GND, __A13_NET_311, __A13_NET_304, __A13_NET_299, __A13_NET_300, __A13_NET_267, CTROR, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U13014(__A13_NET_268, __A13_NET_267, __A13_NET_255, __A13_NET_255, __A13_NET_268, F07A, GND, __A13_NET_255, F07B_n, __A13_NET_257, NHALGA, __A13_1__CKTAL_n, ALGA, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U13015(__A13_NET_297, GNHNC, PSEUDO, __A13_NET_294, PHS2_n, __A13_NET_293, GND, F05B_n, __A13_NET_252, __A13_NET_251, __A13_NET_251, __A13_NET_259, __A13_NET_262, VCC, SIM_RST, SIM_CLK);
    U74HC04 U13016(VFAIL, __A13_NET_252, __A13_NET_260, __A13_1__MVFAIL_n, DBLTEST, __A13_1__CON1, GND, __A13_1__MSCDBL_n, __A13_1__SCADBL, __A13_NET_181, F14B, __A13_1__FILTIN, __A13_NET_178, VCC, SIM_RST, SIM_CLK);
    U74HC27 U13017(__A13_NET_262, __A13_NET_252, F05A_n, __A13_NET_262, NHVFAL, __A13_NET_260, GND, __A13_NET_175, F05A_n, __A13_NET_262, STNDBY_n, __A13_NET_259, NHVFAL, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U13018(__A13_NET_261, __A13_NET_260, STRT1, STRT1, __A13_NET_261, __A13_NET_258, GND, __A13_NET_259, F05A_n, __A13_NET_258, __A13_1__CON3, n2FSFAL, __A13_1__SCADBL, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U13019(__A13_NET_175, __A13_1__DOFILT, SB0_n, __A13_NET_182, __A13_NET_181, __A13_NET_179, GND, __A13_NET_158, FLTOUT, SCAFAL, AGCWAR, __A13_NET_168, __A13_1__SCADBL, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U13020(__A13_1__CON3, __A13_1__CON2, FS10, __A13_1__CON2, __A13_1__CON1, FS09, GND, ALTEST, __A13_NET_169, __A13_NET_170, __A13_NET_182, __A13_NET_171, __A13_NET_169, VCC, SIM_RST, SIM_CLK);
    assign __A13_NET_182 = __A13_NET_182_U13021_2;
    assign __A13_NET_182 = __A13_NET_182_U13021_4;
    assign __A13_NET_266 = __A13_NET_266_U13021_6;
    assign __A13_NET_266 = __A13_NET_266_U13021_8;
    assign __A13_NET_266 = __A13_NET_266_U13021_10;
    assign __A13_NET_266 = __A13_NET_266_U13021_12;
    U74LVC07 U13021(__A13_NET_168, __A13_NET_182_U13021_2, __A13_NET_170, __A13_NET_182_U13021_4, __A13_NET_189, __A13_NET_266_U13021_6, GND, __A13_NET_266_U13021_8, __A13_NET_188, __A13_NET_266_U13021_10, __A13_NET_200, __A13_NET_266_U13021_12, __A13_NET_199, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U13022(__A13_NET_171, SB2_n, __A13_NET_181, __A13_NET_178, __A13_NET_179, __A13_NET_180, GND, __A13_NET_178, F08B, __A13_NET_180, FLTOUT, SCAFAL, __A13_NET_160, VCC, SIM_RST, SIM_CLK);
    U74HC04 U13023(__A13_NET_160, __A13_1__WARN, __A13_1__WARN, __A13_1__CGCWAR, SCAFAL, __A13_1__MSCAFL_n, GND, __A13_1__MWARNF_n, FLTOUT, __A13_1__MOSCAL_n, STRT2, __A13_1__TMPCAU, __A13_NET_166, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U13024(AGCWAR, __A13_NET_158, CCH33, __A13_NET_159, STRT2, OSCALM, GND, __A13_NET_159, CCH33, OSCALM, TEMPIN_n, TMPOUT, __A13_NET_166, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U13025(__A13_NET_162, GOJAM, __A13_NET_167, __A13_NET_161, ALTEST, __A13_NET_162, GND, SBY, __A13_NET_164, __A13_NET_163, __A13_NET_163, T10, __A13_NET_164, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U13026(__A13_NET_162, GOJAM, CT_n, P02_n, P03, __A13_NET_208, GND, __A13_NET_210, T02_n, CA6_n, XB7_n, __A13_NET_167, __A13_1__SBYEXT, VCC, SIM_RST, SIM_CLK);
    U74HC04 U13027(__A13_NET_161, __A13_1__RESTRT, __A13_NET_163, __A13_1__SBYEXT, PIPAFL, __A13_1__MPIPAL_n, GND, __A13_1__SYNC4_n, __A13_NET_207, __A13_1__SYNC14_n, __A13_NET_208, __A13_NET_219, F17A, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U13028(__A13_NET_207, FS01, P02, P03_n, CT_n,  , GND,  , T1P, T2P, T3P, T4P, __A13_NET_206, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U13029(__A13_NET_220, __A13_NET_210, __A13_NET_209, __A13_NET_209, __A13_NET_220, F17B, GND, __A13_NET_219, SB1_n, __A13_NET_213, __A13_1__WATCHP, __A13_1__WATCH, __A13_NET_214, VCC, SIM_RST, SIM_CLK);
    U74HC27 U13030(SB2_n, __A13_NET_209, __A13_NET_304, __A13_NET_302, __A13_NET_300, __A13_NET_301, GND, __A13_NET_291, __A13_NET_304, __A13_NET_292, __A13_NET_300, __A13_1__WATCHP, __A13_NET_219, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b1) U13031(__A13_1__WATCH, __A13_NET_214, __A13_NET_213, __A13_NET_202, OTLNKM, ALTM, GND, __A13_NET_294, __A13_NET_280, __A13_NET_300, __A13_NET_311, __A13_NET_308, __A13_NET_309, VCC, SIM_RST, SIM_CLK);
    U74HC04 U13032(__A13_1__WATCH, __A13_1__MWATCH_n, __A13_NET_303, __A13_NET_304, MLOAD, __A13_NET_299, GND, __A13_NET_302, MREAD, __A13_NET_292, MLDCH, __A13_NET_290, MRDCH, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U13033(__A13_NET_192, T5P, T6P, CDUXP, CDUXM,  , GND,  , CDUYP, CDUYM, CDUZP, CDUZM, __A13_NET_193, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U13034(__A13_NET_187, TRNP, TRNM, SHAFTP, SHAFTM,  , GND,  , PIPXP, PIPXM, PIPYP, PIPYM, __A13_NET_189, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U13035(__A13_NET_188, PIPZP, PIPZM, BMAGXP, BMAGXM,  , GND,  , BMAGYP, BMAGYM, BMAGZP, BMAGZM, __A13_NET_200, VCC, SIM_RST, SIM_CLK);
    assign __A13_NET_266 = __A13_NET_266_U13036_2;
    assign __A13_NET_266 = __A13_NET_266_U13036_4;
    assign __A13_NET_266 = __A13_NET_266_U13036_6;
    assign __A13_NET_303 = __A13_NET_303_U13036_8;
    assign __A13_NET_303 = __A13_NET_303_U13036_10;
    U74LVC07 U13036(__A13_NET_198, __A13_NET_266_U13036_2, __A13_NET_197, __A13_NET_266_U13036_4, __A13_NET_202, __A13_NET_266_U13036_6, GND, __A13_NET_303_U13036_8, __A13_NET_298, __A13_NET_303_U13036_10, __A13_NET_297,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U13037(__A13_NET_304, __A13_NET_290, __A13_NET_300, GOJAM, __A13_NET_276, __A13_NET_280, GND, __A13_NET_308, __A13_NET_309, GOJAM, __A13_NET_306, __A13_NET_289, __A13_NET_300, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U13038(__A13_NET_293, MRDCH, MLDCH, MREAD, MLOAD,  , GND,  , __A13_NET_308, __A13_NET_312, INOTLD, __A13_2__INOTRD, __A13_NET_274, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b0, 1'b1) U13039(__A13_NET_310, __A13_NET_301, __A13_NET_312, __A13_NET_313, __A13_NET_291, INOTLD, GND, __A13_NET_313, __A13_NET_305, INOTLD, __A13_NET_289, __A13_2__INOTRD, __A13_NET_307, VCC, SIM_RST, SIM_CLK);
    U74HC27 U13040(__A13_NET_310, GOJAM, MON_n, __A13_NET_277, ST1_n, __A13_NET_306, GND, __A13_NET_305, T12_n, CT, PHS2_n, __A13_NET_312, __A13_NET_306, VCC, SIM_RST, SIM_CLK);
    U74HC02 U13041(__A13_2__INOTRD, __A13_NET_307, __A13_NET_305, __A13_2__STORE1, ST1_n, __A13_NET_309, GND, ST1_n, __A13_NET_310, FETCH1, __A13_NET_308, __A13_NET_312, MON_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U13042(FETCH0, ST1_n, MON_n, STFET1_n, __A13_2__STORE1, FETCH1, GND, __A13_NET_275, T11_n, __A13_NET_276, CTROR_n, __A13_NET_280, __A13_NET_281, VCC, SIM_RST, SIM_CLK);
    U74HC04 U13043(__A13_NET_305, __A13_NET_277, __A13_2__STORE1, STORE1_n, FETCH0, FETCH0_n, GND, MONpCH, __A13_NET_274, __A13_2__MREQIN, __A13_NET_274, INCSET_n, __A13_NET_286, VCC, SIM_RST, SIM_CLK);
    U74HC27 U13044(FETCH1, __A13_2__STORE1, __A13_NET_281, T12_n, PHS3_n, __A13_NET_288, GND, __A13_NET_287, __A13_NET_285, __A13_NET_288, GOJAM, __A13_NET_275, CHINC, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U13045(__A13_NET_284, __A13_NET_304, MNHNC, __A13_NET_280, CTROR_n,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U13046(__A13_NET_285, __A13_NET_284, __A13_NET_287, __A13_NET_286, T02_n, __A13_NET_285, GND, __A13_NET_287, MONpCH, INKL_n, __A13_2__INOTRD, INOTLD, CHINC_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U13047(INKL_n, INKL, INKL_n, __A13_2__MINKL, T10_n, BKTF_n, GND, CHINC, CHINC_n, __A13_1__FS13_n, FS13,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U13048(__A13_NET_285, T07_n,  ,  ,  ,  , GND,  ,  ,  ,  , RSSB, PHS3_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b1) U14001(__A14_1__ROP_n, S11, S12, __A14_NET_210, T08_n, PHS3_n, GND, __A14_NET_210, __A14_NET_211, __A14_NET_209, __A14_NET_212, __A14_NET_213, __A14_NET_206, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14002(__A14_NET_209, T09, __A14_1__ROP_n, __A14_NET_209, T08, __A14_NET_212, GND, __A14_NET_213, __A14_NET_206, __A14_NET_207, TIMR, __A14_NET_211, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14003(T01_n, __A14_NET_207, __A14_NET_206, __A14_1__IHENV, __A14_NET_219, __A14_1__SETAB_n, GND, SETAB, __A14_1__SETAB_n, __A14_1__SETCD_n, __A14_NET_220, SETCD, __A14_1__SETCD_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14004(TIMR, __A14_NET_207, PHS4_n, __A14_1__ROP_n, T10_n, __A14_NET_208, GND, __A14_NET_214, T05_n, PHS3_n, __A14_1__ROP_n, __A14_NET_205, __A14_NET_218, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U14005(__A14_NET_218, __A14_NET_205, __A14_NET_208, __A14_NET_219, S09, __A14_NET_218, GND, __A14_NET_218, S09_n, __A14_NET_220, __A14_NET_214, __A14_NET_215, __A14_NET_199, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14006(__A14_NET_199, T08, __A14_NET_199, S09, S08, __A14_NET_216, GND, __A14_NET_196, __A14_NET_199, S09, S08_n, __A14_NET_215, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74HC02 U14007(__A14_NET_217, __A14_1__CLEARA, __A14_NET_216, __A14_NET_198, __A14_1__CLEARB, __A14_NET_196, GND, __A14_1__CLEARC, __A14_NET_200, __A14_NET_202, __A14_1__CLEARD, __A14_NET_194, __A14_NET_192, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14008(__A14_NET_217, RESETA, __A14_NET_198, RESETB, __A14_NET_202, RESETC, GND, RESETD, __A14_NET_192, __A14_1__S08A_n, S08, __A14_1__S08A, S08_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U14009(__A14_NET_199, S08, __A14_NET_199, S09_n, S08_n, __A14_NET_194, GND, STBF, GOJAM, __A14_NET_204, __A14_NET_203, __A14_NET_200, S09_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U14010(__A14_1__CLEARA, __A14_1__SETAB_n, __A14_1__S08A_n, __A14_1__CLEARB, __A14_1__SETAB_n, __A14_1__S08A, GND, __A14_1__SETCD_n, __A14_1__S08A_n, __A14_1__CLEARC, __A14_1__SETCD_n, __A14_1__S08A, __A14_1__CLEARD, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U14011(__A14_NET_203, STBF, __A14_1__SBFSET, __A14_NET_204, T07_n, PHS3_n, GND, T02_n, __A14_1__ROP_n, __A14_NET_235, __A14_NET_235, STRGAT, __A14_NET_236, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14012(__A14_NET_203, SBF, __A14_1__ROP_n, __A14_NET_260, S07_n, __A14_2__IL07_n, GND, WEX, __A14_NET_250, WEY, __A14_NET_249, __A14_1__ERAS_n, __A14_1__ERAS, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14013(MNHSBF, MP1, __A14_1__ROP_n, T05_n, DV3764, __A14_NET_280, GND, STRGAT, __A14_NET_236, T08, GOJAM, __A14_NET_279, PHS4_n, VCC, SIM_RST, SIM_CLK);
    assign __A14_1__SBFSET = __A14_1__SBFSET_U14014_2;
    assign __A14_1__SBFSET = __A14_1__SBFSET_U14014_4;
    assign __A14_1__TPGF = __A14_1__TPGF_U14014_6;
    assign __A14_1__TPGF = __A14_1__TPGF_U14014_8;
    assign __A14_1__ERAS = __A14_1__ERAS_U14014_10;
    assign __A14_1__ERAS = __A14_1__ERAS_U14014_12;
    U74LVC07 U14014(__A14_NET_279, __A14_1__SBFSET_U14014_2, __A14_NET_280, __A14_1__SBFSET_U14014_4, __A14_NET_285, __A14_1__TPGF_U14014_6, GND, __A14_1__TPGF_U14014_8, __A14_NET_286, __A14_1__ERAS_U14014_10, __A14_NET_231, __A14_1__ERAS_U14014_12, __A14_NET_226, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U14015(__A14_NET_285, __A14_1__ROP_n, T08_n, DV3764, GOJ1,  , GND,  , GOJAM, TCSAJ3, PHS2_n, MP1, __A14_NET_286, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14016(T02_n, __A14_NET_260, __A14_NET_265, T03, GOJAM, __A14_NET_258, GND, __A14_NET_263, __A14_NET_262, T07, GOJAM, __A14_NET_264, __A14_NET_265, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U14017(__A14_NET_259, __A14_1__ROP_n, T10_n, __A14_NET_265, __A14_NET_259, __A14_NET_258, GND, __A14_NET_264, __A14_NET_263, __A14_NET_262, T01, __A14_NET_261, __A14_NET_253, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U14018(__A14_NET_261, __A14_NET_253, __A14_NET_252, __A14_NET_252, T12_n, PHS3_n, GND, T12A, __A14_NET_261, __A14_NET_257, __A14_NET_251, __A14_NET_255, __A14_NET_250, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14019(__A14_NET_257, TIMR, __A14_NET_257, TIMR, __A14_NET_249, __A14_NET_248, GND, __A14_NET_254, TIMR, T11, __A14_NET_256, __A14_NET_251, __A14_NET_250, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b0, 1'b0) U14020(__A14_NET_249, __A14_NET_248, __A14_NET_276, __A14_NET_256, __A14_NET_254, __A14_NET_270, GND, __A14_NET_256, T10, __A14_NET_255, T05_n, __A14_1__ERAS_n, __A14_NET_275, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14021(__A14_NET_242, __A14_NET_224, __A14_1__ERAS_n, PHS3_n, T03_n, __A14_NET_223, GND, __A14_NET_274, __A14_1__FNERAS_n, T12A, GOJAM, __A14_NET_232, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U14022(__A14_1__FNERAS_n, __A14_NET_275, __A14_NET_274, __A14_NET_271, __A14_1__FNERAS_n, T10_n, GND, __A14_NET_266, __A14_NET_270, __A14_NET_269, T02_n, PHS4_n, __A14_NET_268, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14023(T10_n, __A14_1__FNERAS_n, __A14_1__FNERAS_n, T10_n, PHS3_n, __A14_NET_270, GND, __A14_NET_266, TIMR, __A14_NET_268, __A14_NET_269, __A14_NET_276, PHS4_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14024(TIMR, T01, __A14_NET_222, GOJAM, __A14_1__REDRST, __A14_NET_221, GND, __A14_NET_225, __A14_NET_233, GOJAM, __A14_1__REDRST, __A14_NET_272, __A14_NET_267, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U14025(__A14_NET_267, __A14_NET_272, __A14_NET_271, ZID, __A14_NET_267, STRT2, GND, __A14_1__ERAS_n, T03_n, __A14_NET_234, __A14_NET_234, __A14_NET_232, __A14_NET_242, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U14026(__A14_NET_231, TCSAJ3, S11, S12, INOUT,  , GND,  , CHINC, GOJ1, MP1, MAMU, __A14_NET_226, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b1) U14027(SETEK, STRT2, __A14_NET_242, __A14_NET_224, T06_n, PHS3_n, GND, __A14_NET_223, __A14_NET_221, __A14_NET_222, __A14_NET_237, __A14_NET_225, __A14_NET_233, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14028(__A14_NET_222, __A14_1__REY, __A14_NET_233, __A14_1__REX, __A14_NET_239, SBE, GND, __A14_1__RSTK_n, __A14_NET_269, __A14_1__RSTKY_n, __A14_1__RSTK_n, __A14_1__RSTKX_n, __A14_1__RSTK_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14029(__A14_1__ERAS_n, T03_n, GOJAM, T05, __A14_NET_239, STBE, GND, __A14_1__SBESET, T04_n, __A14_1__ERAS_n, SCAD, __A14_NET_237, PHS4_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U14030(__A14_1__REDRST, __A14_NET_238, T05, __A14_NET_238, __A14_NET_241, __A14_NET_240, GND, __A14_NET_238, T06, __A14_NET_240, T05_n, PHS3_n, __A14_NET_241, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U14031(__A14_NET_239, STBE, __A14_1__SBESET, __A14_NET_247, T05_n, PHS3_n, GND, __A14_1__TPGF, __A14_1__TPGE, TPARG_n, S07, S08, __A14_2__YB0, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14032(SCAD, __A14_1__ERAS_n, S01, S02, S03, XB0, GND, XB1, S01_n, S02, S03, __A14_NET_246, GOJAM, VCC, SIM_RST, SIM_CLK);
    assign __A14_1__TPGE = __A14_1__TPGE_U14033_2;
    assign __A14_1__TPGE = __A14_1__TPGE_U14033_4;
    U74LVC07 U14033(__A14_NET_246, __A14_1__TPGE_U14033_2, __A14_NET_247, __A14_1__TPGE_U14033_4,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U14034(XB0, XB0_n, XB0_n, __A14_2__XB0E, XB1, XB1_n, GND, XB1E, XB1_n, XB2_n, XB2, XB2E, XB2_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14035(S01, S02_n, S01_n, S02_n, S03, XB3, GND, XB4, S01, S02, S03_n, XB2, S03, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14036(XB3, XB3_n, XB3_n, XB3E, XB4, XB4_n, GND, XB4E, XB4_n, XB5_n, XB5, XB5E, XB5_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14037(S01_n, S02, S01, S02_n, S03_n, XB6, GND, XB7, S01_n, S02_n, S03_n, XB5, S03_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14038(XB6, XB6_n, XB6_n, XB6E, XB7, XB7_n, GND, XB7E, XB7_n, YB0_n, __A14_2__YB0, __A14_2__YB0E, YB0_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U14039(__A14_2__YB1, S07_n, S08, __A14_2__YB2, S07, S08_n, GND, S07_n, S08_n, __A14_2__YB3, EB9, S10_n, __A14_NET_287, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14040(__A14_2__YB1, __A14_2__YB1_n, __A14_2__YB1_n, YB1E, __A14_2__YB2, __A14_2__YB2_n, GND, YB2E, __A14_2__YB2_n, __A14_2__YB3_n, __A14_2__YB3, YB3E, __A14_2__YB3_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14041(S04, S05, S04_n, S05, S06, __A14_2__XT1, GND, __A14_2__XT2, S04, S05_n, S06, __A14_2__XT0, S06, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14042(__A14_2__XT0, XT0_n, XT0_n, __A14_2__XT0E, __A14_2__XT1, XT1_n, GND, XT1E, XT1_n, XT2_n, __A14_2__XT2, XT2E, XT2_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14043(S04_n, S05_n, S04, S05, S06_n, __A14_2__XT4, GND, __A14_2__XT5, S04_n, S05, S06_n, __A14_2__XT3, S06, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14044(__A14_2__XT3, XT3_n, XT3_n, XT3E, __A14_2__XT4, XT4_n, GND, XT4E, XT4_n, XT5_n, __A14_2__XT5, XT5E, XT5_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14045(S04, S05_n, S04_n, S05_n, S06_n, __A14_2__XT7, GND, __A14_2__EAD11, S09_n, S10_n, EB11_n, __A14_2__XT6, S06_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14046(__A14_2__XT6, XT6_n, XT6_n, XT6E, __A14_2__XT7, __A14_2__XT7_n, GND, XT7E, __A14_2__XT7_n, __A14_2__EAD09_n, __A14_2__EAD09, __A14_2__EAD10_n, __A14_2__EAD10, VCC, SIM_RST, SIM_CLK);
    U74HC02 U14047(__A14_2__EAD09, __A14_NET_287, S09_n, __A14_NET_306, EB10, S09_n, GND, S10_n, __A14_NET_306, __A14_2__EAD10, __A14_2__YB0, __A14_2__YB3, __A14_2__RILP1, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14048(__A14_2__EAD11, __A14_2__EAD11_n, __A14_2__YT0, YT0_n, YT0_n, __A14_2__YT0E, GND, __A14_2__YT1_n, __A14_2__YT1, YT1E, __A14_2__YT1_n, __A14_2__YT2_n, __A14_2__YT2, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14049(__A14_2__EAD09, __A14_2__EAD10, __A14_2__EAD09_n, __A14_2__EAD10, __A14_2__EAD11, __A14_2__YT1, GND, __A14_2__YT2, __A14_2__EAD09, __A14_2__EAD10_n, __A14_2__EAD11, __A14_2__YT0, __A14_2__EAD11, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14050(__A14_2__YT2_n, YT2E, __A14_2__YT3, __A14_2__YT3_n, __A14_2__YT3_n, YT3E, GND, __A14_2__YT4_n, __A14_2__YT4, YT4E, __A14_2__YT4_n, __A14_2__YT5_n, __A14_2__YT5, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14051(__A14_2__EAD09_n, __A14_2__EAD10_n, __A14_2__EAD09, __A14_2__EAD10, __A14_2__EAD11_n, __A14_2__YT4, GND, __A14_2__YT5, __A14_2__EAD09_n, __A14_2__EAD10, __A14_2__EAD11_n, __A14_2__YT3, __A14_2__EAD11, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14052(__A14_2__YT5_n, YT5E, __A14_2__YT6, __A14_2__YT6_n, __A14_2__YT6_n, YT6E, GND, __A14_2__YT7_n, __A14_2__YT7, YT7E, __A14_2__YT7_n, __A14_NET_288, __A14_NET_292, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14053(__A14_2__EAD09, __A14_2__EAD10_n, __A14_2__EAD09_n, __A14_2__EAD10_n, __A14_2__EAD11_n, __A14_2__YT7, GND, __A14_NET_290, __A14_NET_292, __A14_2__RILP1, __A14_NET_289, __A14_2__YT6, __A14_2__EAD11_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U14054(__A14_NET_292, XB0, XB3, XB5, XB6,  , GND,  , __A14_2__XT0, __A14_2__XT3, __A14_2__XT5, __A14_2__XT6, __A14_NET_289, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14055(__A14_NET_289, __A14_NET_308, __A14_2__RILP1, __A14_2__RILP1_n, __A14_NET_300, __A14_NET_301, GND, __A14_2__ILP_n, __A14_NET_300, __A14_2__ILP, __A14_NET_301, IL01, S01, VCC, SIM_RST, SIM_CLK);
    U74HC27 U14056(__A14_NET_288, __A14_2__RILP1, __A14_NET_288, __A14_2__RILP1_n, __A14_NET_289, __A14_NET_297, GND, __A14_NET_296, __A14_NET_292, __A14_2__RILP1_n, __A14_NET_308, __A14_NET_295, __A14_NET_308, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U14057(__A14_NET_300, __A14_NET_290, __A14_NET_295, __A14_NET_297, __A14_NET_296,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U14058(S01_n, __A14_2__IL01_n, S02, IL02, S02_n, __A14_2__IL02_n, GND, IL03, S03, __A14_2__IL03_n, S03_n, IL04, S04, VCC, SIM_RST, SIM_CLK);
    U74HC04 U14059(S04_n, __A14_2__IL04_n, S05, IL05, S05_n, __A14_2__IL05_n, GND, IL06, S06, __A14_2__IL06_n, S06_n, IL07, S07, VCC, SIM_RST, SIM_CLK);
    U74HC02 U14060(CLROPE, STRT2, __A14_NET_262,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U15001(__A15_NET_168, WL16_n, WFBG_n, __A15_1__FB16, __A15_1__FB16_n, CFBG, GND, __A15_1__FB16_n, RFBG_n, __A15_1__BK16, WL14_n, WFBG_n, __A15_NET_169, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U15002(__A15_NET_168, __A15_NET_167, SUMA16_n, U2BBKG_n, SUMB16_n, __A15_NET_167, GND, __A15_NET_164, SUMA14_n, U2BBKG_n, SUMB14_n, __A15_1__FB16_n, __A15_1__FB16, VCC, SIM_RST, SIM_CLK);
    U74HC04 U15003(__A15_1__BK16, __A15_NET_202, __A15_1__BK16, __A15_NET_203, __A15_NET_163, __A15_NET_204, GND, __A15_NET_199, __A15_NET_175, __A15_NET_212, __A15_NET_151, __A15_NET_205, __A15_NET_162, VCC, SIM_RST, SIM_CLK);
    assign RL16_n = RL16_n_U15004_2;
    assign RL15_n = RL15_n_U15004_4;
    assign RL14_n = RL14_n_U15004_6;
    assign RL13_n = RL13_n_U15004_8;
    assign RL12_n = RL12_n_U15004_10;
    assign RL11_n = RL11_n_U15004_12;
    U74LVC07 U15004(__A15_NET_202, RL16_n_U15004_2, __A15_NET_203, RL15_n_U15004_4, __A15_NET_204, RL14_n_U15004_6, GND, RL13_n_U15004_8, __A15_NET_199, RL12_n_U15004_10, __A15_NET_198, RL11_n_U15004_12, __A15_NET_200, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U15005(__A15_NET_169, __A15_NET_164, SUMA13_n, U2BBKG_n, SUMB13_n, __A15_NET_165, GND, __A15_1__FB13_n, __A15_NET_166, __A15_NET_165, __A15_1__FB13, __A15_1__FB14_n, __A15_1__FB14, VCC, SIM_RST, SIM_CLK);
    U74HC02 U15006(__A15_1__FB14, __A15_1__FB14_n, CFBG, __A15_NET_163, __A15_1__FB14_n, RFBG_n, GND, WL13_n, WFBG_n, __A15_NET_166, __A15_1__FB13_n, CFBG, __A15_1__FB13, VCC, SIM_RST, SIM_CLK);
    U74HC02 U15007(__A15_NET_175, __A15_1__FB13_n, RFBG_n, __A15_NET_174, WL12_n, WFBG_n, GND, __A15_1__FB12_n, CFBG, __A15_1__FB12, __A15_1__FB12_n, RFBG_n, __A15_NET_172, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U15008(SUMA12_n, U2BBKG_n, __A15_NET_174, __A15_NET_176, __A15_1__FB12, __A15_1__FB12_n, GND, __A15_NET_198, RSTRT, __A15_NET_172, __A15_1__RPTA12, __A15_NET_176, SUMB12_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U15009(__A15_NET_171, WFBG_n, WL11_n, __A15_1__FB11, __A15_1__FB11_n, CFBG, GND, __A15_1__FB11_n, RFBG_n, __A15_NET_173, __A15_NET_173, __A15_NET_155, __A15_NET_200, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U15010(SUMA11_n, U2BBKG_n, __A15_NET_171, __A15_NET_170, __A15_1__FB11, __A15_1__FB11_n, GND, __A15_NET_152, SUMA03_n, U2BBKG_n, SUMB03_n, __A15_NET_170, SUMB11_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U15011(__A15_NET_154, WL11_n, WEBG_n, __A15_NET_153, WL03_n, WBBEG_n, GND, EB11_n, CEBG, __A15_1__EB11, REBG_n, EB11_n, __A15_NET_155, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U15012(EB11_n, __A15_NET_152, __A15_NET_154, __A15_NET_153, __A15_1__EB11,  , GND,  , __A15_NET_156, __A15_NET_150, __A15_NET_149, EB10, __A15_1__EB10_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U15013(__A15_1__BBK3, EB11_n, RBBEG_n, __A15_NET_150, WL10_n, WEBG_n, GND, WL02_n, WBBEG_n, __A15_NET_149, __A15_1__EB10_n, CEBG, EB10, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15014(SUMA02_n, U2BBKG_n, SUMA01_n, U2BBKG_n, SUMB01_n, __A15_NET_161, GND, __A15_1__F14, __A15_NET_189, __A15_NET_191, __A15_1__FB14_n, __A15_NET_156, SUMB02_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U15015(__A15_NET_151, REBG_n, __A15_1__EB10_n, __A15_1__BBK2, __A15_1__EB10_n, RBBEG_n, GND, WL09_n, WEBG_n, __A15_NET_159, WL01_n, WBBEG_n, __A15_NET_160, VCC, SIM_RST, SIM_CLK);
    assign RL10_n = RL10_n_U15016_2;
    assign RL09_n = RL09_n_U15016_4;
    assign RL06_n = RL06_n_U15016_6;
    assign __A15_NET_237 = __A15_NET_237_U15016_8;
    assign __A15_NET_237 = __A15_NET_237_U15016_10;
    assign __A15_NET_230 = __A15_NET_230_U15016_12;
    U74LVC07 U15016(__A15_NET_212, RL10_n_U15016_2, __A15_NET_205, RL09_n_U15016_4, __A15_NET_184, RL06_n_U15016_6, GND, __A15_NET_237_U15016_8, __A15_NET_296, __A15_NET_237_U15016_10, __A15_NET_302, __A15_NET_230_U15016_12, __A15_NET_301, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U15017(__A15_1__EB9_n, __A15_NET_161, __A15_NET_159, __A15_NET_160, EB9,  , GND,  , __A15_1__FB14_n, __A15_1__FB16_n, E7_n, __A15_NET_189, __A15_1__F16, VCC, SIM_RST, SIM_CLK);
    U74HC02 U15018(EB9, __A15_1__EB9_n, CEBG, __A15_NET_162, REBG_n, __A15_1__EB9_n, GND, __A15_1__EB9_n, RBBEG_n, __A15_1__BBK1, __A15_1__FB11_n, __A15_NET_189, __A15_NET_158, VCC, SIM_RST, SIM_CLK);
    U74HC04 U15019(S12_n, __A15_NET_189, __A15_1__F11_n, __A15_1__F11, __A15_1__F12_n, __A15_1__F12, GND, __A15_1__F13_n, __A15_1__F13, __A15_1__F14_n, __A15_1__F14, __A15_1__F15_n, __A15_1__F15, VCC, SIM_RST, SIM_CLK);
    U74HC02 U15020(__A15_1__F11_n, __A15_NET_158, __A15_NET_157, __A15_NET_157, S11_n, S12_n, GND, __A15_NET_189, __A15_1__FB12, __A15_1__F12_n, __A15_NET_189, __A15_1__FB13_n, __A15_1__F13, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15021(E5, __A15_1__FB16_n, __A15_1__FB16_n, __A15_NET_192, __A15_NET_189, __A15_1__F15, GND, __A15_NET_192, E7_n, __A15_1__FB14_n, E6, __A15_NET_191, E7_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U15022(__A15_1__F16, __A15_1__F16_n, __A15_NET_252, __A15_NET_224, KRPT, __A15_1__KRPTA_n, GND, __A15_NET_227, __A15_NET_228, __A15_NET_279, __A15_NET_231, __A15_1__PRPOR1, __A15_NET_280, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15023(XB4_n, XT4_n, __A15_1__KRPTA_n, XB0_n, XT5_n, __A15_NET_197, GND, __A15_NET_194, __A15_NET_193, __A15_NET_195, GOJAM, __A15_NET_195, __A15_1__KRPTA_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b0) U15024(__A15_NET_193, RADRPT, __A15_NET_194, __A15_NET_180, HNDRPT, __A15_NET_196, GND, __A15_NET_179, __A15_1__RRPA1_n, __A15_1__RPTAD6, __A15_1__RRPA1_n, __A15_NET_183, __A15_1__RPTA12, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15025(__A15_NET_180, __A15_NET_197, __A15_1__PRPOR1, __A15_NET_193, __A15_1__DNRPTA, __A15_1__PRPOR3, GND, __A15_NET_179, __A15_1__PRPOR2, __A15_1__PRPOR3, __A15_1__PRPOR4, __A15_NET_196, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U15026(__A15_1__PRPOR4, __A15_1__PRPOR1, __A15_1__DNRPTA, __A15_NET_194, __A15_NET_180,  , GND,  , __A15_NET_196, __A15_NET_194, __A15_1__PRPOR1, __A15_1__DNRPTA, __A15_NET_183, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U15027(__A15_NET_184, CAD6, __A15_1__RPTAD6, __A15_NET_185, __A15_NET_183, RUPTOR_n, GND, __A15_NET_185, T10, RUPTOR_n, WOVR_n, OVF_n, __A15_NET_252, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15028(CA3_n, XB1_n, __A15_NET_253, GOJAM, __A15_NET_261, __A15_NET_254, GND, __A15_NET_261, XT0_n, XB4_n, __A15_1__KRPTA_n, __A15_2__T6RPT, ZOUT_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b1) U15029(__A15_NET_253, __A15_2__T6RPT, __A15_NET_254, __A15_NET_258, __A15_NET_260, __A15_NET_256, GND, __A15_NET_220, __A15_NET_219, __A15_NET_218, __A15_NET_223, __A15_NET_225, __A15_NET_222, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15030(CA3_n, XB0_n, __A15_NET_258, GOJAM, __A15_NET_257, __A15_NET_256, GND, __A15_NET_257, XB0_n, XT1_n, __A15_1__KRPTA_n, __A15_NET_260, __A15_NET_224, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15031(CA2_n, XB6_n, __A15_NET_218, GOJAM, __A15_NET_217, __A15_NET_219, GND, __A15_NET_217, XT1_n, XB4_n, __A15_1__KRPTA_n, __A15_NET_220, __A15_NET_224, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15032(CA2_n, XB7_n, __A15_NET_222, GOJAM, __A15_NET_221, __A15_NET_225, GND, __A15_NET_221, XT2_n, XB0_n, __A15_1__KRPTA_n, __A15_NET_223, __A15_NET_224, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b0) U15033(__A15_NET_213, KYRPT1, __A15_NET_214, __A15_NET_235, UPRUPT, __A15_NET_215, GND, DLKPLS, __A15_1__DNRPTA, __A15_NET_233, __A15_NET_254, __A15_NET_258, __A15_NET_229, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U15034(__A15_NET_213, GOJAM, XB4_n, XT2_n, __A15_1__KRPTA_n, __A15_2__KY1RST, GND, __A15_NET_216, KYRPT2, MKRPT, __A15_NET_278, __A15_NET_214, __A15_2__KY1RST, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15035(__A15_NET_216, GOJAM, XT3_n, XB0_n, __A15_1__KRPTA_n, __A15_2__KY2RST, GND, __A15_NET_215, __A15_NET_235, GOJAM, __A15_NET_234, __A15_NET_278, __A15_2__KY2RST, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15036(XT3_n, XB4_n, __A15_NET_233, GOJAM, DRPRST, __A15_1__DNRPTA, GND, DRPRST, XB0_n, XT4_n, __A15_1__KRPTA_n, __A15_NET_234, __A15_1__KRPTA_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U15037(__A15_NET_296, __A15_NET_254, __A15_NET_236, __A15_NET_301, __A15_NET_229, __A15_NET_236, GND, __A15_NET_227, __A15_NET_222, __A15_NET_226, __A15_NET_279, __A15_NET_216, __A15_NET_282, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15038(__A15_NET_232, __A15_NET_281, __A15_NET_254, __A15_NET_218, __A15_NET_256, __A15_NET_236, GND, __A15_NET_298, __A15_NET_282, __A15_NET_281, __A15_1__PRPOR4, __A15_NET_302, __A15_1__PRPOR3, VCC, SIM_RST, SIM_CLK);
    assign __A15_NET_230 = __A15_NET_230_U15039_2;
    assign RL03_n = RL03_n_U15039_4;
    assign RL04_n = RL04_n_U15039_6;
    assign RL05_n = RL05_n_U15039_8;
    assign RL02_n = RL02_n_U15039_10;
    assign RL01_n = RL01_n_U15039_12;
    U74LVC07 U15039(__A15_NET_298, __A15_NET_230_U15039_2, __A15_NET_304, RL03_n_U15039_4, __A15_NET_307, RL04_n_U15039_6, GND, RL05_n_U15039_8, __A15_NET_308, RL02_n_U15039_10, __A15_NET_306, RL01_n_U15039_12, __A15_NET_305, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15040(__A15_NET_254, __A15_NET_219, __A15_NET_227, __A15_NET_213, __A15_NET_225, __A15_NET_232, GND, __A15_NET_231, __A15_NET_227, __A15_NET_214, __A15_NET_225, __A15_NET_228, __A15_NET_256, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U15041(__A15_NET_246, __A15_NET_232, __A15_NET_226, __A15_NET_282, __A15_NET_281,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U15042(__A15_NET_279, __A15_NET_235, __A15_NET_279, __A15_NET_215, __A15_NET_278, __A15_NET_280, GND, __A15_NET_304, __A15_2__RPTAD3, __A15_1__BBK3, CAD3, __A15_NET_281, __A15_NET_278, VCC, SIM_RST, SIM_CLK);
    U74HC02 U15043(__A15_1__PRPOR2, __A15_1__PRPOR1, __A15_NET_233, __A15_2__RPTAD3, __A15_1__RRPA1_n, __A15_NET_237, GND, __A15_1__RRPA1_n, __A15_NET_230, __A15_2__RPTAD4, __A15_2__RPTAD4, CAD4, __A15_NET_307, VCC, SIM_RST, SIM_CLK);
    U74HC04 U15044(RRPA, __A15_1__RRPA1_n, STRGAT, __A15_NET_277, __A15_1__F11, __A15_NET_276, GND, __A15_NET_291, __A15_1__F11_n, __A15_NET_290, S10, __A15_NET_289, S10_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U15045(__A15_NET_308, __A15_2__RPTAD5, CAD5,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U15046(CAD2, __A15_1__BBK2, CAD1, __A15_1__BBK1, RB1F, __A15_NET_305, GND, STR412, __A15_NET_277, __A15_NET_290, __A15_NET_276, __A15_NET_306, R6, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15047(__A15_NET_277, __A15_NET_289, __A15_NET_277, __A15_NET_290, __A15_NET_291, STR210, GND, STR19, __A15_NET_277, __A15_NET_289, __A15_NET_291, STR311, __A15_NET_276, VCC, SIM_RST, SIM_CLK);
    U74HC02 U15048(__A15_NET_288, __A15_1__F16, __A15_1__F15, __A15_NET_286, __A15_1__F16, __A15_1__F15_n, GND, __A15_1__F15, __A15_1__F16_n, __A15_NET_245, __A15_2__NE036_n, __A15_1__F12, __A15_2__036L, VCC, SIM_RST, SIM_CLK);
    U74HC04 U15049(__A15_NET_288, __A15_NET_294, __A15_1__F14_n, __A15_NET_295, __A15_1__F13_n, __A15_NET_293, GND, __A15_NET_292, __A15_1__F13, __A15_NET_284, __A15_1__F14, __A15_NET_285, __A15_NET_286, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15050(__A15_NET_294, __A15_NET_295, __A15_NET_294, __A15_NET_295, __A15_NET_292, __A15_2__NE01, GND, __A15_2__NE02, __A15_NET_294, __A15_NET_284, __A15_NET_293, __A15_2__NE00, __A15_NET_293, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15051(__A15_NET_294, __A15_NET_284, __A15_NET_285, __A15_NET_295, __A15_NET_293, __A15_2__NE04, GND, __A15_2__NE05, __A15_NET_285, __A15_NET_295, __A15_NET_292, __A15_2__NE03, __A15_NET_292, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15052(__A15_NET_285, __A15_NET_284, __A15_NET_285, __A15_NET_284, __A15_NET_292, __A15_2__NE07, GND, __A15_2__NE10, __A15_NET_287, __A15_NET_295, __A15_NET_293, __A15_2__NE06, __A15_NET_293, VCC, SIM_RST, SIM_CLK);
    U74HC04 U15053(__A15_NET_245, __A15_NET_287, __A15_NET_263, STR14, __A15_2__NE012_n, ROPER, GND, LOMOD, __A15_NET_273, STR58, __A15_NET_274, ROPES, __A15_2__NE345_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15054(__A15_2__NE00, __A15_2__NE03, __A15_2__NE00, __A15_2__NE01, __A15_2__NE02, __A15_2__NE012_n, GND, __A15_2__NE147_n, __A15_2__NE01, __A15_2__NE04, __A15_2__NE07, __A15_2__NE036_n, __A15_2__NE06, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15055(__A15_2__NE04, __A15_2__NE03, __A15_2__NE02, __A15_2__NE05, __A15_2__NE10, __A15_2__NE2510_n, GND, __A15_2__NE6710_n, __A15_2__NE06, __A15_2__NE07, __A15_2__NE10, __A15_2__NE345_n, __A15_2__NE05, VCC, SIM_RST, SIM_CLK);
    U74HC02 U15056(__A15_2__147H, __A15_2__NE147_n, __A15_1__F12_n, __A15_2__2510L, __A15_2__NE2510_n, __A15_1__F12, GND, __A15_2__NE036_n, __A15_1__F12_n, __A15_2__036H, __A15_2__NE147_n, __A15_1__F12, __A15_2__147L, VCC, SIM_RST, SIM_CLK);
    U74HC02 U15057(__A15_2__2510H, __A15_2__NE2510_n, __A15_1__F12_n, __A15_NET_263, __A15_2__036L, __A15_2__147H, GND, __A15_2__2510L, __A15_2__036H, __A15_NET_274, __A15_2__147L, __A15_2__2510H, __A15_NET_255, VCC, SIM_RST, SIM_CLK);
    U74HC27 U15058(__A15_2__036L, __A15_2__147L, __A15_2__147H, __A15_2__2510H, __A15_2__2510L, __A15_NET_270, GND,  ,  ,  ,  , __A15_NET_273, __A15_2__036H, VCC, SIM_RST, SIM_CLK);
    U74HC04 U15059(__A15_NET_270, HIMOD, __A15_NET_255, STR912, __A15_2__NE6710_n, ROPET, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U15060(__A15_2__RPTAD5, __A15_1__RRPA1_n, __A15_NET_246,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16001(__A16_NET_117, CHWL01_n, __A16_1__WCH05_n, __A16_NET_118, __A16_NET_117, __A16_NET_116, GND, __A16_NET_118, __A16_1__CCH05, __A16_NET_116, __A16_NET_118, __A16_1__RCH05_n, __A16_NET_122, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16002(__A16_NET_118, __A16_1__RCpXpP, __A16_NET_119, __A16_1__RCpZpR, __A16_NET_108, __A16_1__RCmXmP, GND, __A16_1__RCmZmR, __A16_NET_113, __A16_1__RCmXpP, __A16_NET_133, __A16_1__RCmZpR, __A16_NET_124, VCC, SIM_RST, SIM_CLK);
    U74HC27 U16003(__A16_NET_111, __A16_NET_122, __A16_NET_129, __A16_NET_112, CH3202, __A16_NET_196, GND, __A16_NET_193, __A16_NET_123, __A16_NET_132, CH3203, __A16_NET_195, CH3201, VCC, SIM_RST, SIM_CLK);
    assign __A16_1__CHOR01_n = __A16_1__CHOR01_n_U16004_2;
    assign __A16_1__CHOR02_n = __A16_1__CHOR02_n_U16004_4;
    assign __A16_1__CHOR03_n = __A16_1__CHOR03_n_U16004_6;
    assign __A16_1__CHOR04_n = __A16_1__CHOR04_n_U16004_8;
    assign __A16_1__CHOR05_n = __A16_1__CHOR05_n_U16004_10;
    assign __A16_1__CHOR06_n = __A16_1__CHOR06_n_U16004_12;
    U74LVC07 U16004(__A16_NET_195, __A16_1__CHOR01_n_U16004_2, __A16_NET_196, __A16_1__CHOR02_n_U16004_4, __A16_NET_193, __A16_1__CHOR03_n_U16004_6, GND, __A16_1__CHOR04_n_U16004_8, __A16_NET_194, __A16_1__CHOR05_n_U16004_10, __A16_NET_199, __A16_1__CHOR06_n_U16004_12, __A16_NET_200, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16005(__A16_NET_121, CHWL01_n, __A16_1__WCH06_n, __A16_NET_119, __A16_NET_121, __A16_NET_120, GND, __A16_NET_119, __A16_1__CCH06, __A16_NET_120, __A16_NET_119, __A16_1__RCH06_n, __A16_NET_111, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16006(__A16_NET_110, CHWL02_n, __A16_1__WCH05_n, __A16_NET_108, __A16_NET_110, __A16_NET_109, GND, __A16_NET_108, __A16_1__CCH05, __A16_NET_109, __A16_NET_108, __A16_1__RCH05_n, __A16_NET_112, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16007(__A16_NET_115, CHWL02_n, __A16_1__WCH06_n, __A16_NET_113, __A16_NET_115, __A16_NET_114, GND, __A16_NET_113, __A16_NET_128, __A16_NET_114, __A16_NET_113, __A16_1__RCH06_n, __A16_NET_129, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16008(__A16_NET_135, CHWL03_n, __A16_1__WCH05_n, __A16_NET_133, __A16_NET_135, __A16_NET_134, GND, __A16_NET_133, __A16_1__CCH05, __A16_NET_134, __A16_NET_133, __A16_1__RCH05_n, __A16_NET_132, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16009(__A16_NET_131, CHWL03_n, __A16_1__WCH06_n, __A16_NET_124, __A16_NET_131, __A16_NET_130, GND, __A16_NET_124, __A16_1__CCH06, __A16_NET_130, __A16_NET_124, __A16_1__RCH06_n, __A16_NET_123, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16010(__A16_NET_127, CHWL04_n, __A16_1__WCH05_n, __A16_NET_125, __A16_NET_127, __A16_NET_126, GND, __A16_NET_125, __A16_1__CCH05, __A16_NET_126, __A16_NET_125, __A16_1__RCH05_n, __A16_NET_172, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16011(__A16_NET_125, __A16_1__RCpXmP, __A16_NET_169, __A16_1__RCpZmR, __A16_NET_163, __A16_1__RCpXpY, GND, __A16_1__RCpYpR, __A16_NET_161, __A16_1__RCmXmY, __A16_NET_186, __A16_1__RCmYmR, __A16_NET_191, VCC, SIM_RST, SIM_CLK);
    U74HC27 U16012(__A16_NET_177, __A16_NET_172, __A16_NET_167, __A16_NET_162, CH3205, __A16_NET_199, GND, __A16_NET_200, __A16_NET_182, __A16_NET_188, CH3206, __A16_NET_194, CH3204, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16013(__A16_NET_171, CHWL04_n, __A16_1__WCH06_n, __A16_NET_169, __A16_NET_171, __A16_NET_170, GND, __A16_NET_169, __A16_1__CCH06, __A16_NET_170, __A16_NET_169, __A16_1__RCH06_n, __A16_NET_177, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16014(__A16_NET_174, CHWL05_n, __A16_1__WCH05_n, __A16_NET_163, __A16_NET_174, __A16_NET_168, GND, __A16_NET_163, __A16_1__CCH05, __A16_NET_168, __A16_NET_163, __A16_1__RCH05_n, __A16_NET_162, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16015(__A16_NET_160, CHWL05_n, __A16_1__WCH06_n, __A16_NET_161, __A16_NET_160, __A16_NET_159, GND, __A16_NET_161, __A16_1__CCH06, __A16_NET_159, __A16_NET_161, __A16_1__RCH06_n, __A16_NET_167, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16016(__A16_NET_190, CHWL06_n, __A16_1__WCH05_n, __A16_NET_186, __A16_NET_190, __A16_NET_189, GND, __A16_NET_186, __A16_1__CCH05, __A16_NET_189, __A16_NET_186, __A16_1__RCH05_n, __A16_NET_188, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16017(__A16_NET_187, CHWL06_n, __A16_1__WCH06_n, __A16_NET_191, __A16_NET_187, __A16_NET_192, GND, __A16_NET_191, __A16_1__CCH06, __A16_NET_192, __A16_NET_191, __A16_1__RCH06_n, __A16_NET_182, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16018(__A16_NET_179, CHWL07_n, __A16_1__WCH05_n, __A16_NET_185, __A16_NET_179, __A16_NET_178, GND, __A16_NET_185, __A16_1__CCH05, __A16_NET_178, __A16_NET_185, __A16_1__RCH05_n, __A16_NET_184, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16019(__A16_NET_185, __A16_1__RCmXpY, __A16_NET_181, __A16_1__RCmYpR, __A16_NET_157, __A16_1__RCpXmY, GND, __A16_1__RCpYmR, __A16_NET_151, __A16_1__WCH05_n, __A16_NET_138, __A16_1__WCH06_n, __A16_NET_140, VCC, SIM_RST, SIM_CLK);
    U74HC27 U16020(__A16_NET_153, __A16_NET_184, __A16_NET_150, __A16_NET_156, CH3208, __A16_NET_198, GND, __A16_NET_138, WCHG_n, XT0_n, XB5_n, __A16_NET_197, CH3207, VCC, SIM_RST, SIM_CLK);
    assign __A16_1__CHOR07_n = __A16_1__CHOR07_n_U16021_2;
    assign __A16_1__CHOR08_n = __A16_1__CHOR08_n_U16021_4;
    assign __A16_2__CHOR01_n = __A16_2__CHOR01_n_U16021_6;
    assign __A16_2__CHOR02_n = __A16_2__CHOR02_n_U16021_8;
    assign __A16_2__CHOR03_n = __A16_2__CHOR03_n_U16021_10;
    assign __A16_2__CHOR04_n = __A16_2__CHOR04_n_U16021_12;
    U74LVC07 U16021(__A16_NET_197, __A16_1__CHOR07_n_U16021_2, __A16_NET_198, __A16_1__CHOR08_n_U16021_4, __A16_NET_270, __A16_2__CHOR01_n_U16021_6, GND, __A16_2__CHOR02_n_U16021_8, __A16_NET_267, __A16_2__CHOR03_n_U16021_10, __A16_NET_266, __A16_2__CHOR04_n_U16021_12, __A16_NET_268, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16022(__A16_NET_183, CHWL07_n, __A16_1__WCH06_n, __A16_NET_181, __A16_NET_183, __A16_NET_180, GND, __A16_NET_181, __A16_1__CCH06, __A16_NET_180, __A16_NET_181, __A16_1__RCH06_n, __A16_NET_153, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16023(__A16_NET_152, CHWL08_n, __A16_1__WCH05_n, __A16_NET_157, __A16_NET_152, __A16_NET_158, GND, __A16_NET_157, __A16_1__CCH05, __A16_NET_158, __A16_NET_157, __A16_1__RCH05_n, __A16_NET_156, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16024(__A16_NET_155, CHWL08_n, __A16_1__WCH06_n, __A16_NET_151, __A16_NET_155, __A16_NET_154, GND, __A16_NET_151, __A16_1__CCH06, __A16_NET_154, __A16_NET_151, __A16_1__RCH06_n, __A16_NET_150, VCC, SIM_RST, SIM_CLK);
    U74HC27 U16025(WCHG_n, XT0_n, CCHG_n, XT0_n, XB5_n, __A16_NET_139, GND, __A16_NET_146, CCHG_n, XT0_n, XB6_n, __A16_NET_140, XB6_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16026(__A16_NET_136, __A16_1__CCH05, __A16_NET_137, __A16_1__RCH05_n, __A16_NET_144, __A16_1__RCH06_n, GND, __A16_1__CCH06, __A16_NET_145, __A16_1__TVCNAB, __A16_NET_147, __A16_1__OT1207, __A16_NET_142, VCC, SIM_RST, SIM_CLK);
    U74HC02 U16027(__A16_NET_136, __A16_NET_139, GOJAM, __A16_NET_137, XT0_n, XB5_n, GND, XT0_n, XB6_n, __A16_NET_144, __A16_NET_146, GOJAM, __A16_NET_145, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16028(__A16_NET_149, CHWL08_n, __A16_1__WCH12_n, __A16_NET_147, __A16_NET_149, __A16_NET_148, GND, __A16_NET_147, __A16_1__CCH12, __A16_NET_148, __A16_1__RCH12_n, __A16_NET_147, __A16_1__CH1208, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16029(__A16_NET_143, __A16_1__WCH12_n, CHWL07_n, __A16_NET_142, __A16_NET_143, __A16_NET_141, GND, __A16_NET_142, __A16_1__CCH12, __A16_NET_141, __A16_1__RCH12_n, __A16_NET_142, __A16_1__CH1207, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16030(__A16_NET_141, __A16_1__OT1207_n, __A16_NET_274, __A16_2__ZOPCDU, __A16_NET_273, __A16_2__ZOPCDU, GND, __A16_2__ENEROP, __A16_NET_233, __A16_2__COMACT, __A16_NET_236, __A16_2__STARON, __A16_NET_225, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16031(__A16_NET_276, CHWL01_n, __A16_1__WCH12_n, __A16_NET_274, __A16_NET_276, __A16_NET_275, GND, __A16_NET_274, __A16_1__CCH12, __A16_NET_275, __A16_NET_274, __A16_1__RCH12_n, __A16_NET_272, VCC, SIM_RST, SIM_CLK);
    U74HC27 U16032(__A16_NET_272, __A16_NET_271, __A16_NET_235, __A16_NET_234, CH1502, __A16_NET_267, GND, __A16_NET_266, __A16_NET_244, __A16_NET_243, CH1503, __A16_NET_270, CH1501, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16033(__A16_NET_277, CHWL01_n, WCH11_n, __A16_NET_273, __A16_NET_277, __A16_NET_269, GND, __A16_NET_273, CCH11, __A16_NET_269, __A16_NET_273, RCH11_n, __A16_NET_271, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16034(__A16_NET_278, CHWL02_n, __A16_1__WCH12_n, __A16_NET_233, __A16_NET_278, __A16_NET_279, GND, __A16_NET_233, __A16_1__CCH12, __A16_NET_279, __A16_NET_233, __A16_1__RCH12_n, __A16_NET_235, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16035(__A16_NET_232, CHWL02_n, WCH11_n, __A16_NET_236, __A16_NET_232, __A16_NET_231, GND, __A16_NET_236, CCH11, __A16_NET_231, __A16_NET_236, RCH11_n, __A16_NET_234, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16036(__A16_NET_227, CHWL03_n, __A16_1__WCH12_n, __A16_NET_225, __A16_NET_227, __A16_NET_226, GND, __A16_NET_225, __A16_1__CCH12, __A16_NET_226, __A16_NET_225, __A16_1__RCH12_n, __A16_NET_244, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16037(__A16_NET_230, CHWL03_n, WCH11_n, __A16_NET_228, __A16_NET_230, __A16_NET_229, GND, __A16_NET_228, CCH11, __A16_NET_229, __A16_NET_228, RCH11_n, __A16_NET_243, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16038(__A16_NET_228, __A16_2__UPLACT, __A16_NET_248, __A16_2__COARSE, __A16_NET_245, TMPOUT, GND, __A16_2__ZIMCDU, __A16_NET_239, __A16_2__ENERIM, __A16_NET_204, __A16_2__S4BTAK, __A16_NET_220, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16039(__A16_NET_242, CHWL04_n, __A16_1__WCH12_n, __A16_NET_248, __A16_NET_242, __A16_NET_249, GND, __A16_NET_248, __A16_1__CCH12, __A16_NET_249, __A16_NET_248, __A16_1__RCH12_n, __A16_NET_238, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16040(__A16_NET_247, CHWL04_n, WCH11_n, __A16_NET_245, __A16_NET_247, __A16_NET_246, GND, __A16_NET_245, CCH11, __A16_NET_246, __A16_NET_245, RCH11_n, __A16_NET_237, VCC, SIM_RST, SIM_CLK);
    U74HC27 U16041(__A16_NET_238, __A16_NET_237, __A16_NET_207, __A16_NET_213, CH0705, __A16_NET_281, GND, __A16_NET_280, __A16_NET_206, __A16_NET_205, CH0706, __A16_NET_268, CH1504, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16042(__A16_NET_241, CHWL05_n, __A16_1__WCH12_n, __A16_NET_239, __A16_NET_241, __A16_NET_240, GND, __A16_NET_239, __A16_1__CCH12, __A16_NET_240, __A16_NET_239, __A16_1__RCH12_n, __A16_NET_207, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16043(__A16_NET_210, CHWL05_n, WCH11_n, __A16_NET_208, __A16_NET_210, __A16_NET_209, GND, __A16_NET_208, CCH11, __A16_NET_209, __A16_NET_208, RCH11_n, __A16_NET_213, VCC, SIM_RST, SIM_CLK);
    assign __A16_2__CHOR05_n = __A16_2__CHOR05_n_U16044_2;
    assign __A16_2__CHOR06_n = __A16_2__CHOR06_n_U16044_4;
    assign __A16_2__CHOR07_n = __A16_2__CHOR07_n_U16044_6;
    U74LVC07 U16044(__A16_NET_281, __A16_2__CHOR05_n_U16044_2, __A16_NET_280, __A16_2__CHOR06_n_U16044_4, __A16_NET_265, __A16_2__CHOR07_n_U16044_6, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16045(__A16_NET_212, CHWL06_n, __A16_1__WCH12_n, __A16_NET_204, __A16_NET_212, __A16_NET_211, GND, __A16_NET_204, __A16_1__CCH12, __A16_NET_211, __A16_NET_204, __A16_1__RCH12_n, __A16_NET_206, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16046(__A16_NET_203, CHWL06_n, WCH11_n, __A16_NET_201, __A16_NET_203, __A16_NET_202, GND, __A16_NET_201, CCH11, __A16_NET_202, __A16_NET_201, RCH11_n, __A16_NET_205, VCC, SIM_RST, SIM_CLK);
    U74HC02 U16047(__A16_2__KYRLS, __A16_NET_208, FLASH, __A16_2__VNFLSH, __A16_NET_201, FLASH_n, GND, __A16_NET_264, FLASH, __A16_2__OPEROR, __A16_NET_261, GOJAM, __A16_NET_262, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16048(__A16_NET_221, CHWL09_n, __A16_1__WCH12_n, __A16_NET_220, __A16_NET_221, __A16_NET_219, GND, __A16_NET_220, __A16_1__CCH12, __A16_NET_219, __A16_NET_220, __A16_1__RCH12_n, __A16_2__CH1209, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16049(__A16_NET_224, CHWL10_n, __A16_1__WCH12_n, __A16_NET_223, __A16_NET_224, __A16_NET_222, GND, __A16_NET_223, __A16_1__CCH12, __A16_NET_222, __A16_NET_223, __A16_1__RCH12_n, __A16_2__CH1210, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16050(__A16_NET_223, __A16_2__ZEROPT, __A16_NET_215, __A16_2__DISDAC, __A16_NET_255, __A16_2__MROLGT, GND, __A16_2__S4BSEQ, __A16_NET_257, __A16_2__S4BOFF, __A16_NET_250, __A16_1__WCH12_n, __A16_NET_253, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16051(__A16_NET_216, CHWL11_n, __A16_1__WCH12_n, __A16_NET_215, __A16_NET_216, __A16_NET_214, GND, __A16_NET_215, __A16_1__CCH12, __A16_NET_214, __A16_NET_215, __A16_1__RCH12_n, __A16_2__CH1211, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16052(__A16_NET_218, CHWL07_n, WCH11_n, __A16_NET_264, __A16_NET_218, __A16_NET_217, GND, __A16_NET_264, CCH11, __A16_NET_217, __A16_NET_264, RCH11_n, __A16_NET_263, VCC, SIM_RST, SIM_CLK);
    U74HC27 U16053(__A16_1__CH1207, __A16_NET_263, WCHG_n, XB2_n, XT1_n, __A16_NET_253, GND, __A16_NET_261, CCHG_n, XB2_n, XT1_n, __A16_NET_265, CH0707, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16054(__A16_NET_256, CHWL12_n, __A16_1__WCH12_n, __A16_NET_255, __A16_NET_256, __A16_NET_254, GND, __A16_NET_255, __A16_1__CCH12, __A16_NET_254, __A16_NET_255, __A16_1__RCH12_n, __A16_2__CH1212, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16055(__A16_NET_259, CHWL13_n, __A16_1__WCH12_n, __A16_NET_257, __A16_NET_259, __A16_NET_258, GND, __A16_NET_257, __A16_1__CCH12, __A16_NET_258, __A16_NET_257, __A16_1__RCH12_n, CH1213, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16056(__A16_NET_252, CHWL14_n, __A16_1__WCH12_n, __A16_NET_250, __A16_NET_252, __A16_NET_251, GND, __A16_NET_250, __A16_1__CCH12, __A16_NET_251, __A16_NET_250, __A16_1__RCH12_n, CH1214, VCC, SIM_RST, SIM_CLK);
    U74HC04 U16057(__A16_NET_262, __A16_1__CCH12, __A16_NET_260, __A16_1__RCH12_n,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U16058(__A16_NET_260, XT1_n, XB2_n,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U17001(__A17_NET_226, IN3301, __A17_1__RCH33_n, __A17_NET_227, XB3_n, XT3_n, GND, ULLTHR, __A17_1__RCH30_n, __A17_NET_224, XB0_n, XT3_n, __A17_NET_251, VCC, SIM_RST, SIM_CLK);
    U74HC04 U17002(__A17_NET_227, __A17_1__RCH33_n, __A17_NET_251, __A17_1__RCH30_n, __A17_NET_225, __A17_1__RCH31_n, GND, __A17_1__RCH32_n, __A17_NET_215, __A17_1__F04B_n, F04B, __A17_2__RLYB01, __A17_NET_346, VCC, SIM_RST, SIM_CLK);
    assign __A17_1__CHOR01_n = __A17_1__CHOR01_n_U17004_2;
    assign __A17_1__CHOR02_n = __A17_1__CHOR02_n_U17004_4;
    assign __A17_1__CHOR03_n = __A17_1__CHOR03_n_U17004_6;
    assign __A17_1__CHOR04_n = __A17_1__CHOR04_n_U17004_8;
    assign __A17_1__CHOR05_n = __A17_1__CHOR05_n_U17004_10;
    assign __A17_1__CHOR06_n = __A17_1__CHOR06_n_U17004_12;
    U74LVC07 U17004(__A17_NET_273, __A17_1__CHOR01_n_U17004_2, __A17_NET_272, __A17_1__CHOR02_n_U17004_4, __A17_NET_275, __A17_1__CHOR03_n_U17004_6, GND, __A17_1__CHOR04_n_U17004_8, __A17_NET_274, __A17_1__CHOR05_n_U17004_10, __A17_NET_268, __A17_1__CHOR06_n_U17004_12, __A17_NET_266, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17005(__A17_NET_230, MANpP, __A17_1__RCH31_n, __A17_NET_225, XB1_n, XT3_n, GND, SMSEPR, __A17_1__RCH30_n, __A17_NET_228, RRPONA, __A17_1__RCH33_n, __A17_NET_229, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17006(__A17_NET_219, MANmP, __A17_1__RCH31_n, __A17_NET_218, RRRLSC, __A17_1__RCH33_n, GND, MANpY, __A17_1__RCH31_n, __A17_NET_216, SPSRDY, __A17_1__RCH30_n, __A17_NET_217, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17007(__A17_NET_226, __A17_NET_224, __A17_NET_229, __A17_NET_228, __A17_NET_219, __A17_NET_272, GND, __A17_NET_275, __A17_NET_218, __A17_NET_217, __A17_NET_216, __A17_NET_273, __A17_NET_230, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17008(__A17_NET_222, S4BSAB, __A17_1__RCH30_n, __A17_NET_223, ZEROP, __A17_1__RCH33_n, GND, MANmY, __A17_1__RCH31_n, __A17_NET_221, LFTOFF, __A17_1__RCH30_n, __A17_NET_241, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17009(__A17_NET_223, __A17_NET_222, __A17_NET_220, __A17_NET_241, __A17_NET_240, __A17_NET_268, GND, __A17_NET_266, __A17_NET_239, __A17_NET_238, __A17_NET_245, __A17_NET_274, __A17_NET_221, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17010(__A17_NET_220, OPMSW2, __A17_1__RCH33_n, __A17_NET_240, MANpR, __A17_1__RCH31_n, GND, GUIREL, __A17_1__RCH30_n, __A17_NET_238, OPMSW3, __A17_1__RCH33_n, __A17_NET_239, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17011(__A17_NET_245, MANmR, __A17_1__RCH31_n, __A17_NET_243, OPCDFL, __A17_1__RCH30_n, GND, STRPRS, __A17_1__RCH33_n, __A17_NET_244, TRANpX, __A17_1__RCH31_n, __A17_NET_242, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17012(__A17_NET_244, __A17_NET_243, __A17_NET_234, __A17_NET_233, __A17_NET_232, __A17_NET_271, GND, __A17_NET_269, __A17_NET_231, __A17_NET_237, __A17_NET_236, __A17_NET_267, __A17_NET_242, VCC, SIM_RST, SIM_CLK);
    assign __A17_1__CHOR07_n = __A17_1__CHOR07_n_U17013_2;
    assign __A17_1__CHOR08_n = __A17_1__CHOR08_n_U17013_4;
    assign __A17_1__CHOR09_n = __A17_1__CHOR09_n_U17013_6;
    assign __A17_1__CHOR10_n = __A17_1__CHOR10_n_U17013_8;
    assign __A17_1__CHOR11_n = __A17_1__CHOR11_n_U17013_10;
    assign __A17_1__CHOR12_n = __A17_1__CHOR12_n_U17013_12;
    U74LVC07 U17013(__A17_NET_267, __A17_1__CHOR07_n_U17013_2, __A17_NET_271, __A17_1__CHOR08_n_U17013_4, __A17_NET_269, __A17_1__CHOR09_n_U17013_6, GND, __A17_1__CHOR10_n_U17013_8, __A17_NET_270, __A17_1__CHOR11_n_U17013_10, __A17_NET_282, __A17_1__CHOR12_n_U17013_12, __A17_NET_281, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17014(__A17_NET_233, IN3008, __A17_1__RCH30_n, __A17_NET_234, LVDAGD, __A17_1__RCH33_n, GND, TRANmX, __A17_1__RCH31_n, __A17_NET_232, IMUOPR, __A17_1__RCH30_n, __A17_NET_237, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17015(__A17_NET_231, LRRLSC, __A17_1__RCH33_n, __A17_NET_236, TRANpY, __A17_1__RCH31_n, GND, CTLSAT, __A17_1__RCH30_n, __A17_NET_235, TRANmY, __A17_1__RCH31_n, __A17_NET_200, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17016(CH3310, __A17_NET_235, __A17_NET_199, __A17_NET_198, __A17_NET_197, __A17_NET_282, GND, __A17_NET_281, __A17_NET_205, __A17_NET_204, __A17_NET_203, __A17_NET_270, __A17_NET_200, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17017(__A17_NET_198, IMUCAG, __A17_1__RCH30_n, __A17_NET_199, LEMATT, __A17_1__RCH32_n, GND, TRANpZ, __A17_1__RCH31_n, __A17_NET_197, CDUFAL, __A17_1__RCH30_n, __A17_NET_204, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17018(__A17_NET_205, IN3212, __A17_1__RCH32_n, __A17_NET_203, TRANmZ, __A17_1__RCH31_n, GND, IMUFAL, __A17_1__RCH30_n, __A17_NET_201, IN3213, __A17_1__RCH32_n, __A17_NET_202, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17019(__A17_NET_202, __A17_NET_201, __A17_NET_190, __A17_NET_191, __A17_NET_196, __A17_NET_283, GND, __A17_NET_284, __A17_NET_195, __A17_NET_193, __A17_NET_194, __A17_NET_285, __A17_NET_192, VCC, SIM_RST, SIM_CLK);
    assign __A17_1__CHOR13_n = __A17_1__CHOR13_n_U17020_2;
    assign __A17_1__CHOR14_n = __A17_1__CHOR14_n_U17020_4;
    assign __A17_1__CHOR16_n = __A17_1__CHOR16_n_U17020_6;
    assign __A17_NET_207 = __A17_NET_207_U17020_8;
    assign __A17_NET_207 = __A17_NET_207_U17020_10;
    assign __A17_NET_254 = __A17_NET_254_U17020_12;
    U74LVC07 U17020(__A17_NET_285, __A17_1__CHOR13_n_U17020_2, __A17_NET_283, __A17_1__CHOR14_n_U17020_4, __A17_NET_284, __A17_1__CHOR16_n_U17020_6, GND, __A17_NET_207_U17020_8, __A17_NET_277, __A17_NET_207_U17020_10, __A17_NET_276, __A17_NET_254_U17020_12, __A17_NET_280, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17021(__A17_NET_192, HOLFUN, __A17_1__RCH31_n, __A17_NET_191, ISSTOR, __A17_1__RCH30_n, GND, IN3214, __A17_1__RCH32_n, __A17_NET_190, FREFUN, __A17_1__RCH31_n, __A17_NET_196, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17022(__A17_NET_193, TEMPIN, __A17_1__RCH30_n, __A17_NET_195, IN3216, __A17_1__RCH32_n, GND, GCAPCL, __A17_1__RCH31_n, __A17_NET_194, XB2_n, XT3_n, __A17_NET_215, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17023(MANpP, MANmP, MANmY, MANpR, MANmR, __A17_NET_276, GND, __A17_NET_212, __A17_NET_213, __A17_NET_207, F05A_n, __A17_NET_277, MANpY, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U17024(__A17_NET_210, CHWL12_n, WCH13_n, __A17_NET_213, __A17_NET_210, __A17_NET_214, GND, __A17_NET_212, __A17_NET_211, __A17_NET_209, __A17_1__F04B_n, FS05_n, __A17_1__FO5D, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17025(__A17_NET_213, GOJAM, __A17_NET_209, __A17_NET_207, __A17_1__FO5D, __A17_NET_211, GND, __A17_NET_280, TRANpX, TRANmX, TRANpY, __A17_NET_214, __A17_1__TRP31A, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U17026(__A17_1__TRP31A, __A17_NET_209, F05B_n, __A17_NET_255, __A17_NET_257, __A17_NET_256, GND, CHWL13_n, WCH13_n, __A17_NET_208, __A17_NET_255, F05B_n, __A17_1__TRP31B, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17027(TRANmY, TRANpZ, __A17_NET_258, __A17_NET_254, F05A_n, __A17_NET_257, GND, __A17_NET_256, __A17_NET_255, __A17_NET_254, __A17_1__FO5D, __A17_NET_278, TRANmZ, VCC, SIM_RST, SIM_CLK);
    assign __A17_NET_254 = __A17_NET_254_U17028_2;
    assign __A17_NET_265 = __A17_NET_265_U17028_4;
    assign __A17_NET_265 = __A17_NET_265_U17028_6;
    assign __A17_NET_265 = __A17_NET_265_U17028_8;
    assign __A17_2__CHOR01_n = __A17_2__CHOR01_n_U17028_10;
    assign __A17_2__CHOR07_n = __A17_2__CHOR07_n_U17028_12;
    U74LVC07 U17028(__A17_NET_278, __A17_NET_254_U17028_2, __A17_NET_264, __A17_NET_265_U17028_4, __A17_NET_262, __A17_NET_265_U17028_6, GND, __A17_NET_265_U17028_8, __A17_NET_261, __A17_2__CHOR01_n_U17028_10, __A17_NET_342, __A17_2__CHOR07_n_U17028_12, __A17_NET_356, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17029(__A17_NET_258, GOJAM, MNIMpR, MNIMmR, TRST9, __A17_NET_262, GND, __A17_NET_261, TRST10, PCHGOF, ROLGOF, __A17_NET_259, __A17_1__TRP31B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17030(__A17_NET_258, __A17_NET_208, __A17_NET_259, CH3201, MNIMpP, __A17_1__RCH32_n, GND, MNIMmP, __A17_1__RCH32_n, CH3202, MNIMpY, __A17_1__RCH32_n, CH3203, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17031(CH3204, MNIMmY, __A17_1__RCH32_n, CH3205, MNIMpR, __A17_1__RCH32_n, GND, MNIMmR, __A17_1__RCH32_n, CH3206, TRST9, __A17_1__RCH32_n, CH3207, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U17032(CH3208, TRST10, __A17_1__RCH32_n, __A17_1__CH3209, PCHGOF, __A17_1__RCH32_n, GND, ROLGOF, __A17_1__RCH32_n, __A17_1__CH3210, __A17_NET_250, __A17_NET_249, __A17_NET_248, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U17033(__A17_NET_264, MNIMpP, MNIMmP, MNIMpY, MNIMmY,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U17034(WCHG_n, XT1_n, __A17_NET_252, __A17_NET_265, F05A_n, __A17_NET_250, GND, __A17_NET_249, __A17_NET_248, __A17_1__FO5D, __A17_NET_265, __A17_NET_312, XB1_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U17035(__A17_1__TRP32, __A17_NET_248, F05B_n, __A17_NET_247, CHWL14_n, WCH13_n, GND, __A17_NET_247, __A17_NET_246, __A17_NET_252, __A17_NET_253, TPOR_n, __A17_1__HNDRPT, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17036(__A17_NET_252, GOJAM, __A17_1__TRP31A, __A17_1__TRP31B, __A17_1__TRP32, __A17_NET_253, GND, __A17_NET_342, CH1301, __A17_NET_341, CH1401, __A17_NET_246, __A17_1__TRP32, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17037(__A17_1__CH3313, PIPAFL, __A17_1__RCH33_n, __A17_1__CH3314, AGCWAR, __A17_1__RCH33_n, GND, OSCALM, __A17_1__RCH33_n, __A17_1__CH3316, CHWL01_n, __A17_2__WCH10_n, __A17_NET_344, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17038(__A17_NET_346, __A17_NET_344, __A17_NET_345, __A17_NET_345, __A17_NET_346, __A17_2__CCH10, GND, __A17_NET_346, __A17_2__RCH10_n, __A17_NET_341, CHWL02_n, __A17_2__WCH10_n, __A17_NET_343, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17039(__A17_NET_350, __A17_NET_343, __A17_NET_349, __A17_NET_349, __A17_NET_350, __A17_2__CCH10, GND, __A17_NET_350, __A17_2__RCH10_n, __A17_NET_348, CHWL03_n, __A17_2__WCH10_n, __A17_NET_331, VCC, SIM_RST, SIM_CLK);
    U74HC04 U17040(__A17_NET_350, __A17_2__RLYB02, __A17_NET_332, __A17_2__RLYB03, __A17_NET_339, __A17_2__RLYB04, GND, __A17_2__RLYB05, __A17_NET_336, __A17_2__RLYB06, __A17_NET_369, __A17_2__RLYB07, __A17_NET_368, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17041(CH1302, __A17_NET_348, CH1303, __A17_NET_327, CH1403, __A17_NET_326, GND, __A17_NET_333, CH1304, __A17_NET_340, CH1404, __A17_NET_347, CH1402, VCC, SIM_RST, SIM_CLK);
    assign __A17_2__CHOR02_n = __A17_2__CHOR02_n_U17042_2;
    assign __A17_2__CHOR03_n = __A17_2__CHOR03_n_U17042_4;
    assign __A17_2__CHOR04_n = __A17_2__CHOR04_n_U17042_6;
    assign __A17_2__CHOR05_n = __A17_2__CHOR05_n_U17042_8;
    assign __A17_2__CHOR06_n = __A17_2__CHOR06_n_U17042_10;
    assign __A17_2__CHOR08_n = __A17_2__CHOR08_n_U17042_12;
    U74LVC07 U17042(__A17_NET_347, __A17_2__CHOR02_n_U17042_2, __A17_NET_326, __A17_2__CHOR03_n_U17042_4, __A17_NET_333, __A17_2__CHOR04_n_U17042_6, GND, __A17_2__CHOR05_n_U17042_8, __A17_NET_363, __A17_2__CHOR06_n_U17042_10, __A17_NET_371, __A17_2__CHOR08_n_U17042_12, __A17_NET_360, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17043(__A17_NET_332, __A17_NET_331, __A17_NET_330, __A17_NET_330, __A17_NET_332, __A17_2__CCH10, GND, __A17_NET_332, __A17_2__RCH10_n, __A17_NET_327, CHWL04_n, __A17_2__WCH10_n, __A17_NET_328, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17044(__A17_NET_339, __A17_NET_328, __A17_NET_329, __A17_NET_329, __A17_NET_339, __A17_2__CCH10, GND, __A17_NET_339, __A17_2__RCH10_n, __A17_NET_340, CHWL05_n, __A17_2__WCH10_n, __A17_NET_337, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17045(__A17_NET_336, __A17_NET_337, __A17_NET_334, __A17_NET_334, __A17_NET_336, __A17_2__CCH10, GND, __A17_NET_336, __A17_2__RCH10_n, __A17_NET_365, CHWL06_n, __A17_2__WCH10_n, __A17_NET_361, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17046(CH1305, __A17_NET_365, CH1306, __A17_NET_370, CH1406, __A17_NET_371, GND,  ,  ,  ,  , __A17_NET_363, CH1405, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17047(__A17_NET_369, __A17_NET_361, __A17_NET_364, __A17_NET_364, __A17_NET_369, __A17_2__CCH10, GND, __A17_NET_369, __A17_2__RCH10_n, __A17_NET_370, CHWL07_n, __A17_2__WCH10_n, __A17_NET_366, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17048(__A17_NET_368, __A17_NET_366, __A17_NET_367, __A17_NET_367, __A17_NET_368, __A17_2__CCH10, GND, __A17_NET_368, __A17_2__RCH10_n, __A17_NET_355, CHWL08_n, __A17_2__WCH10_n, __A17_NET_351, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17049(CH1307, __A17_NET_355, CH1308, __A17_NET_354, CH1408, __A17_NET_360, GND, __A17_NET_303, CH1309, __A17_NET_302, CH1409, __A17_NET_356, CH1407, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17050(__A17_NET_353, __A17_NET_351, __A17_NET_352, __A17_NET_352, __A17_NET_353, __A17_2__CCH10, GND, __A17_NET_353, __A17_2__RCH10_n, __A17_NET_354, CHWL09_n, __A17_2__WCH10_n, __A17_NET_359, VCC, SIM_RST, SIM_CLK);
    U74HC04 U17051(__A17_NET_353, __A17_2__RLYB08, __A17_NET_358, __A17_2__RLYB09, __A17_NET_300, __A17_2__RLYB10, GND, __A17_2__RLYB11, __A17_NET_306, __A17_2__RYWD12, __A17_NET_287, __A17_2__RYWD13, __A17_NET_296, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17052(__A17_NET_358, __A17_NET_359, __A17_NET_357, __A17_NET_357, __A17_NET_358, __A17_2__CCH10, GND, __A17_NET_358, __A17_2__RCH10_n, __A17_NET_302, CHWL10_n, __A17_2__WCH10_n, __A17_NET_299, VCC, SIM_RST, SIM_CLK);
    assign __A17_2__CHOR09_n = __A17_2__CHOR09_n_U17053_2;
    assign __A17_2__CHOR10_n = __A17_2__CHOR10_n_U17053_4;
    assign __A17_2__CHOR11_n = __A17_2__CHOR11_n_U17053_6;
    assign __A17_2__CHOR12_n = __A17_2__CHOR12_n_U17053_8;
    assign __A17_2__CHOR13_n = __A17_2__CHOR13_n_U17053_10;
    assign __A17_2__CHOR14_n = __A17_2__CHOR14_n_U17053_12;
    U74LVC07 U17053(__A17_NET_303, __A17_2__CHOR09_n_U17053_2, __A17_NET_307, __A17_2__CHOR10_n_U17053_4, __A17_NET_289, __A17_2__CHOR11_n_U17053_6, GND, __A17_2__CHOR12_n_U17053_8, __A17_NET_288, __A17_2__CHOR13_n_U17053_10, __A17_NET_294, __A17_2__CHOR14_n_U17053_12, __A17_NET_316, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17054(__A17_NET_300, __A17_NET_299, __A17_NET_298, __A17_NET_298, __A17_NET_300, __A17_2__CCH10, GND, __A17_NET_300, __A17_2__RCH10_n, __A17_NET_301, CHWL11_n, __A17_2__WCH10_n, __A17_NET_305, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17055(CH1310, __A17_NET_301, CH1311, __A17_NET_290, CH1411, __A17_NET_289, GND, __A17_NET_288, CH3312, __A17_NET_286, CH1412, __A17_NET_307, CH1410, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17056(__A17_NET_306, __A17_NET_305, __A17_NET_304, __A17_NET_304, __A17_NET_306, __A17_2__CCH10, GND, __A17_NET_306, __A17_2__RCH10_n, __A17_NET_290, CHWL12_n, __A17_2__WCH10_n, __A17_NET_292, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17057(__A17_NET_287, __A17_NET_292, __A17_NET_291, __A17_NET_291, __A17_NET_287, __A17_2__CCH10, GND, __A17_NET_287, __A17_2__RCH10_n, __A17_NET_286, CHWL13_n, __A17_2__WCH10_n, __A17_NET_295, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17058(__A17_NET_296, __A17_NET_295, __A17_NET_297, __A17_NET_297, __A17_NET_296, __A17_2__CCH10, GND, __A17_NET_296, __A17_2__RCH10_n, __A17_NET_293, CHWL14_n, __A17_2__WCH10_n, __A17_NET_318, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17059(__A17_NET_320, __A17_NET_318, __A17_NET_319, __A17_NET_319, __A17_NET_320, __A17_2__CCH10, GND, __A17_NET_320, __A17_2__RCH10_n, __A17_NET_317, CHWL16_n, __A17_2__WCH10_n, __A17_NET_324, VCC, SIM_RST, SIM_CLK);
    U74HC04 U17060(__A17_NET_320, __A17_2__RYWD14, __A17_NET_323, __A17_2__RYWD16, __A17_NET_311, __A17_2__WCH10_n, GND, __A17_2__CCH10, __A17_NET_310, WCH11_n, __A17_NET_312, CCH11, __A17_NET_313, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17061(__A17_NET_323, __A17_NET_324, __A17_NET_325, __A17_NET_325, __A17_NET_323, __A17_2__CCH10, GND, __A17_NET_323, __A17_2__RCH10_n, __A17_NET_321, __A17_NET_309, GOJAM, __A17_NET_310, VCC, SIM_RST, SIM_CLK);
    assign __A17_2__CHOR16_n = __A17_2__CHOR16_n_U17062_2;
    U74LVC07 U17062(__A17_NET_322, __A17_2__CHOR16_n_U17062_2,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U17063(CH1213, __A17_NET_293, CH1214, __A17_NET_317, CH1414, __A17_NET_316, GND, __A17_NET_322, CH1316, __A17_NET_321, CH1416, __A17_NET_294, CH1413, VCC, SIM_RST, SIM_CLK);
    U74HC27 U17064(WCHG_n, XB0_n, CCHG_n, XT1_n, XB0_n, __A17_NET_309, GND, __A17_NET_314, CCHG_n, XT1_n, XB1_n, __A17_NET_311, XT1_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U17065(__A17_NET_308, XT1_n, XB0_n, __A17_NET_313, __A17_NET_314, GOJAM, GND, XT1_n, XB1_n, __A17_NET_315,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC04 U17066(__A17_NET_308, __A17_2__RCH10_n, __A17_NET_315, RCH11_n,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U18001(__A18_NET_126, MKEY1, __A18_NET_125, __A18_NET_125, __A18_NET_126, __A18_NET_112, GND, __A18_NET_126, __A18_1__RCH15_n, CH1501, MKEY2, __A18_NET_98, __A18_NET_97, VCC, SIM_RST, SIM_CLK);
    U74HC04 U18002(__A18_NET_126, __A18_NET_92, __A18_NET_97, __A18_NET_93, __A18_NET_101, __A18_NET_91, GND, __A18_NET_94, __A18_NET_99, __A18_NET_95, __A18_NET_89, __A18_NET_105, MAINRS, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U18003(__A18_NET_98, __A18_NET_97, __A18_NET_112, CH1502, __A18_NET_97, __A18_1__RCH15_n, GND, MKEY3, __A18_NET_96, __A18_NET_101, __A18_NET_101, __A18_NET_112, __A18_NET_96, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18004(CH1503, __A18_NET_101, __A18_1__RCH15_n, __A18_NET_99, MKEY4, __A18_NET_100, GND, __A18_NET_99, __A18_NET_112, __A18_NET_100, __A18_NET_99, __A18_1__RCH15_n, CH1504, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18005(__A18_NET_89, MKEY5, __A18_NET_90, __A18_NET_90, __A18_NET_89, __A18_NET_112, GND, __A18_NET_89, __A18_1__RCH15_n, __A18_1__CH1505, __A18_NET_94, __A18_NET_95, __A18_NET_185, VCC, SIM_RST, SIM_CLK);
    U74HC27 U18006(__A18_NET_92, __A18_NET_93, __A18_NET_109, __A18_NET_111, __A18_1__F09D, __A18_NET_108, GND, KYRPT1, TPOR_n, __A18_NET_109, F09B_n, __A18_NET_184, __A18_NET_91, VCC, SIM_RST, SIM_CLK);
    assign __A18_NET_111 = __A18_NET_111_U18007_2;
    assign __A18_NET_111 = __A18_NET_111_U18007_4;
    assign __A18_NET_153 = __A18_NET_153_U18007_6;
    assign __A18_NET_153 = __A18_NET_153_U18007_8;
    assign __A18_2__CNTOF9 = __A18_2__CNTOF9_U18007_10;
    assign __A18_2__CNTOF9 = __A18_2__CNTOF9_U18007_12;
    U74LVC07 U18007(__A18_NET_184, __A18_NET_111_U18007_2, __A18_NET_185, __A18_NET_111_U18007_4, __A18_NET_186, __A18_NET_153_U18007_6, GND, __A18_NET_153_U18007_8, __A18_NET_190, __A18_2__CNTOF9_U18007_10, __A18_NET_198, __A18_2__CNTOF9_U18007_12, __A18_NET_199, VCC, SIM_RST, SIM_CLK);
    U74HC04 U18008(__A18_NET_105, __A18_NET_112, __A18_NET_113, __A18_1__RCH15_n, __A18_NET_111, __A18_NET_102, GND, __A18_NET_155, NAVRST, __A18_NET_157, __A18_NET_155, __A18_1__RCH16_n, __A18_NET_154, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U18009( ,  ,  , __A18_NET_113, XT1_n, XB5_n, GND, __A18_NET_110, __A18_NET_108, __A18_NET_109, T05, T11, TPOR_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U18010(__A18_NET_110, __A18_1__F09A_n, __A18_NET_111, __A18_NET_112, __A18_NET_114,  , GND,  , __A18_1__F09A_n, __A18_NET_153, __A18_NET_157, __A18_NET_180, __A18_NET_152, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18011(__A18_NET_116, __A18_NET_102, __A18_NET_105, __A18_NET_114, __A18_NET_116, __A18_NET_115, GND, __A18_NET_114, KYRPT1, __A18_NET_115, XT1_n, XB6_n, __A18_NET_154, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U18012(__A18_NET_104, NKEY1, __A18_NET_103, __A18_NET_103, __A18_NET_104, __A18_NET_157, GND, __A18_NET_104, __A18_1__RCH16_n, __A18_1__CH1601, NKEY2, __A18_NET_107, __A18_NET_106, VCC, SIM_RST, SIM_CLK);
    U74HC04 U18013(__A18_NET_104, __A18_NET_147, __A18_NET_106, __A18_NET_148, __A18_NET_158, __A18_NET_149, GND, __A18_NET_150, __A18_NET_162, __A18_NET_151, __A18_NET_160, __A18_NET_176, __A18_NET_153, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U18014(__A18_NET_107, __A18_NET_106, __A18_NET_157, __A18_1__CH1602, __A18_NET_106, __A18_1__RCH16_n, GND, NKEY3, __A18_NET_159, __A18_NET_158, __A18_NET_158, __A18_NET_157, __A18_NET_159, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18015(__A18_1__CH1603, __A18_NET_158, __A18_1__RCH16_n, __A18_NET_162, NKEY4, __A18_NET_156, GND, __A18_NET_162, __A18_NET_157, __A18_NET_156, __A18_NET_162, __A18_1__RCH16_n, __A18_1__CH1604, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18016(__A18_NET_160, NKEY5, __A18_NET_161, __A18_NET_161, __A18_NET_160, __A18_NET_157, GND, __A18_NET_160, __A18_1__RCH16_n, __A18_1__CH1605, __A18_NET_150, __A18_NET_151, __A18_NET_190, VCC, SIM_RST, SIM_CLK);
    U74HC27 U18017(__A18_NET_147, __A18_NET_148, __A18_NET_175, __A18_NET_153, __A18_1__F09D, __A18_NET_174, GND, KYRPT2, TPOR_n, __A18_NET_175, F09B_n, __A18_NET_186, __A18_NET_149, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U18018(__A18_NET_175, __A18_NET_152, __A18_NET_174, __A18_NET_172, __A18_NET_176, __A18_NET_155, GND, __A18_NET_172, __A18_NET_173, __A18_NET_180, __A18_NET_180, KYRPT2, __A18_NET_173, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18019(__A18_NET_177, WCH13_n, CHWL11_n, __A18_NET_178, __A18_NET_177, __A18_NET_179, GND, __A18_NET_178, CCH13, __A18_NET_179, __A18_NET_178, RCH13_n, CH1311, VCC, SIM_RST, SIM_CLK);
    U74HC04 U18020(SBYBUT, __A18_NET_170, F17A, __A18_1__F17A_n, F17B, __A18_1__F17B_n, GND, STNDBY_n, __A18_1__STNDBY, SBY, STNDBY_n, __A18_1__SBYLIT, __A18_NET_120, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18021(__A18_NET_166, __A18_1__F17A_n, __A18_NET_170, __A18_NET_164, __A18_NET_166, __A18_NET_165, GND, __A18_NET_164, __A18_NET_170, __A18_NET_165, __A18_1__F17B_n, __A18_NET_164, __A18_NET_167, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U18022(__A18_NET_168, __A18_NET_167, __A18_NET_169, __A18_NET_169, __A18_NET_168, __A18_NET_170, GND, __A18_NET_141, __A18_NET_143, __A18_NET_142, __A18_NET_142, __A18_NET_168, __A18_NET_143, VCC, SIM_RST, SIM_CLK);
    U74HC27 U18023(__A18_NET_168, STOP, __A18_2__ACTV_n, RADRPT, __A18_NET_242, __A18_NET_216, GND, __A18_2__ADVCNT, F10A_n, __A18_NET_231, SB2_n, __A18_NET_141, __A18_NET_178, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18024(__A18_NET_144, __A18_NET_143, __A18_NET_168, __A18_NET_140, __A18_NET_143, __A18_1__STNDBY, GND, __A18_NET_140, __A18_NET_144, __A18_1__STNDBY, __A18_1__STNDBY, ALTEST, __A18_NET_120, VCC, SIM_RST, SIM_CLK);
    U74HC04 U18025(MRKRST, __A18_NET_138, __A18_NET_138, __A18_NET_121, __A18_NET_122, __A18_NET_119, GND, __A18_NET_118, __A18_NET_139, __A18_NET_136, __A18_NET_131, __A18_1__F08B_n, F08B, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U18026(__A18_NET_122, MARK, __A18_NET_123, __A18_NET_123, __A18_NET_122, __A18_NET_121, GND, MRKREJ, __A18_NET_117, __A18_NET_139, __A18_NET_139, __A18_NET_121, __A18_NET_117, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U18027(__A18_1__CH1606, __A18_NET_122, __A18_1__RCH16_n, __A18_1__CH1607, __A18_NET_139, __A18_1__RCH16_n, GND, __A18_NET_119, __A18_NET_118, __A18_NET_131, __A18_NET_128, __A18_NET_129, __A18_NET_127, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U18028(__A18_NET_128, __A18_1__F09A_n, __A18_NET_131, __A18_NET_121, __A18_NET_134,  , GND,  , __A18_NET_258, RADRPT, __A18_2__ADVCNT, __A18_NET_262, __A18_NET_261, VCC, SIM_RST, SIM_CLK);
    U74HC27 U18029(TPOR_n, __A18_NET_127, __A18_NET_127, __A18_NET_131, __A18_1__F09D, __A18_NET_129, GND,  ,  ,  ,  , MKRPT, F09B_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18030(__A18_NET_137, __A18_NET_136, __A18_NET_138, __A18_NET_134, __A18_NET_137, __A18_NET_124, GND, __A18_NET_134, MKRPT, __A18_NET_124, __A18_NET_146, FS09_n, __A18_1__F09D, VCC, SIM_RST, SIM_CLK);
    U74HC04 U18031(__A18_1__F08B_n, __A18_NET_146, __A18_NET_237, __A18_NET_208, __A18_NET_194, __A18_NET_207, GND, __A18_NET_193, __A18_NET_192, __A18_NET_195, __A18_NET_191, __A18_NET_220, __A18_2__CNTOF9, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18032(__A18_NET_238, CHWL04_n, WCH13_n, __A18_2__ACTV_n, __A18_NET_238, __A18_NET_216, GND, RCH13_n, __A18_2__ACTV_n, CH1304, CHWL03_n, WCH13_n, __A18_NET_236, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18033(__A18_NET_237, __A18_NET_236, __A18_NET_194, __A18_NET_194, __A18_NET_237, __A18_NET_242, GND, RCH13_n, __A18_NET_237, CH1303, CHWL02_n, WCH13_n, __A18_NET_241, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18034(__A18_NET_240, __A18_NET_241, __A18_NET_196, __A18_NET_196, __A18_NET_240, __A18_NET_242, GND, RCH13_n, __A18_NET_240, CH1302, CHWL01_n, WCH13_n, __A18_NET_230, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18035(__A18_NET_229, __A18_NET_230, __A18_NET_221, __A18_NET_221, __A18_NET_229, __A18_NET_242, GND, RCH13_n, __A18_NET_229, CH1301, F10A_n, SB0_n, __A18_2__F10AS0, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18036(__A18_NET_231, __A18_2__F10AS0, __A18_NET_228, __A18_NET_228, __A18_NET_231, __A18_2__ACTV_n, GND, __A18_NET_262, __A18_NET_259, __A18_NET_232, __A18_NET_261, __A18_NET_259, __A18_NET_260, VCC, SIM_RST, SIM_CLK);
    U74HC27 U18037(__A18_NET_261, __A18_2__ADVCNT, __A18_NET_260, RADRPT, __A18_NET_261, __A18_NET_258, GND, __A18_NET_268, __A18_NET_266, __A18_NET_258, __A18_NET_267, __A18_NET_262, __A18_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC02 U18038(__A18_NET_259, __A18_NET_260, __A18_NET_262, __A18_NET_257, __A18_NET_270, __A18_NET_266, GND, __A18_NET_268, __A18_NET_263, __A18_NET_267, __A18_NET_266, __A18_NET_263, __A18_NET_270, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U18039(__A18_NET_266, __A18_NET_257, RADRPT, __A18_NET_258, __A18_NET_268,  , GND,  , __A18_NET_249, RADRPT, __A18_NET_257, __A18_NET_246, __A18_NET_247, VCC, SIM_RST, SIM_CLK);
    U74HC02 U18040(__A18_NET_263, __A18_NET_270, __A18_NET_268, __A18_NET_249, __A18_NET_244, __A18_NET_247, GND, __A18_NET_246, __A18_NET_243, __A18_NET_245, __A18_NET_247, __A18_NET_243, __A18_NET_244, VCC, SIM_RST, SIM_CLK);
    U74HC27 U18041(__A18_NET_247, __A18_NET_257, __A18_NET_251, __A18_NET_249, __A18_NET_250, __A18_NET_252, GND, __A18_NET_199, __A18_NET_263, __A18_NET_260, F10A, __A18_NET_246, __A18_NET_245, VCC, SIM_RST, SIM_CLK);
    U74HC02 U18042(__A18_NET_243, __A18_NET_244, __A18_NET_246, __A18_NET_248, __A18_NET_200, __A18_NET_251, GND, __A18_NET_252, __A18_NET_269, __A18_NET_250, __A18_NET_251, __A18_NET_269, __A18_NET_200, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U18043(__A18_NET_251, __A18_NET_248, RADRPT, __A18_NET_249, __A18_NET_252,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U18044(__A18_NET_269, __A18_NET_200, __A18_NET_252, __A18_NET_198, __A18_NET_200, __A18_NET_243, GND, __A18_2__ADVCNT, __A18_NET_201, __A18_NET_202, __A18_NET_196, __A18_NET_221, __A18_NET_197, VCC, SIM_RST, SIM_CLK);
    U74HC27 U18045(__A18_NET_202, __A18_2__CNTOF9, __A18_NET_208, __A18_NET_202, F5BSB2_n, __A18_NET_192, GND, __A18_NET_191, F5BSB2_n, __A18_NET_202, __A18_NET_207, __A18_NET_201, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74HC27 U18046(__A18_NET_196, __A18_NET_229, __A18_NET_193, __A18_NET_221, __A18_NET_240, __A18_2__RRRARA, GND, __A18_2__LRXVEL, __A18_NET_221, __A18_NET_196, __A18_NET_195, __A18_2__RRRANG, __A18_NET_193, VCC, SIM_RST, SIM_CLK);
    U74HC27 U18047(__A18_NET_195, __A18_NET_229, __A18_NET_195, __A18_NET_240, __A18_NET_221, __A18_2__LRZVEL, GND, __A18_2__LRRANG, __A18_NET_195, __A18_NET_240, __A18_NET_229, __A18_2__LRYVEL, __A18_NET_196, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U18048(__A18_NET_219, __A18_NET_220, GTSET_n, __A18_NET_217, __A18_NET_219, __A18_NET_218, GND, F5ASB2_n, __A18_NET_217, __A18_NET_225, __A18_NET_225, __A18_NET_226, __A18_NET_224, VCC, SIM_RST, SIM_CLK);
    U74HC27 U18049(__A18_NET_217, RADRPT, __A18_NET_224, F09B, GOJAM, __A18_NET_226, GND, RADRPT, __A18_NET_223, __A18_NET_224, GTRST_n, __A18_NET_218, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74HC04 U18050(TPOR_n, __A18_2__HERB, __A18_2__HERB, __A18_NET_223, __A18_NET_209, __A18_NET_203, GND, __A18_NET_205, RRIN1, __A18_NET_204, RRIN0, __A18_NET_206, LRIN1, VCC, SIM_RST, SIM_CLK);
    U74HC02 U18051(__A18_NET_209, __A18_NET_197, __A18_NET_208, RNRADP, __A18_NET_210, __A18_NET_211, GND, __A18_NET_213, __A18_NET_214, RNRADM,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U18052(__A18_NET_203, __A18_NET_205, __A18_NET_203, __A18_NET_204, __A18_NET_212, __A18_NET_213, GND, __A18_NET_211, __A18_NET_207, __A18_NET_206, __A18_NET_212, __A18_NET_210, __A18_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC04 U18053(LRIN0, __A18_NET_215, __A18_NET_216, __A18_NET_212, F09A, __A18_1__F09A_n, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U18054(__A18_NET_207, __A18_NET_215,  ,  ,  ,  , GND,  ,  ,  ,  , __A18_NET_214, __A18_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U19001(__A19_NET_210, CA6_n, CXB0_n, __A19_NET_209, SHINC_n, T06_n, GND, __A19_NET_209, __A19_NET_208, __A19_1__SH3MS_n, __A19_1__SH3MS_n, CSG, __A19_NET_208, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1) U19002(__A19_NET_210, __A19_NET_215, __A19_NET_214, __A19_NET_223, __A19_NET_211, __A19_1__ALTSNC, GND, __A19_NET_234, __A19_NET_236, __A19_1__OTLNK0, __A19_NET_232, __A19_1__F5ASB0_n, __A19_1__F5ASB0, VCC, SIM_RST, SIM_CLK);
    U74HC27 U19003(BR1, __A19_1__SH3MS_n, __A19_NET_215, __A19_1__SH3MS_n, BR1_n, __A19_NET_226, GND, __A19_NET_229, __A19_NET_228, CCH14, __A19_NET_218, __A19_NET_214, __A19_NET_215, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19004(__A19_NET_213, CHWL02_n, WCH14_n, __A19_NET_225, __A19_NET_213, __A19_NET_224, GND, __A19_NET_225, CCH14, __A19_NET_224, RCH14_n, __A19_NET_225, CH1402, VCC, SIM_RST, SIM_CLK);
    U74HC02 U19005(__A19_1__ALT0, __A19_NET_223, __A19_NET_224, __A19_1__ALT1, __A19_NET_224, __A19_NET_230, GND, __A19_NET_223, __A19_NET_225, __A19_1__ALRT0, __A19_NET_225, __A19_NET_230, __A19_1__ALRT1, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U19006(__A19_NET_230, __A19_NET_226, __A19_NET_222, __A19_NET_227, WCH14_n, CHWL03_n, GND, __A19_NET_227, __A19_NET_229, __A19_NET_228, __A19_NET_229, __A19_NET_218, __A19_NET_221, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19007(CH1403, RCH14_n, __A19_NET_221, __A19_NET_220, __A19_NET_216, __A19_NET_231, GND, __A19_NET_228, GTSET_n, __A19_NET_216, F5ASB2_n, __A19_NET_220, __A19_NET_222, VCC, SIM_RST, SIM_CLK);
    U74HC27 U19008(__A19_NET_220, GOJAM, __A19_NET_219, GTSET, GOJAM, __A19_NET_218, GND, __A19_NET_211, __A19_NET_217, __A19_NET_218, __A19_NET_231, __A19_NET_231, GTONE, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U19009(__A19_NET_219, __A19_NET_222, __A19_NET_218, ALTM, __A19_1__F5ASB0_n, __A19_NET_219, GND, __A19_NET_218, __A19_NET_217, __A19_NET_212, __A19_NET_212, GTONE, __A19_NET_217, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U19010(__A19_NET_239, CHWL01_n, WCH14_n, __A19_NET_240, __A19_NET_239, __A19_NET_245, GND, GTSET_n, __A19_NET_240, __A19_NET_243, __A19_NET_243, __A19_NET_242, __A19_NET_241, VCC, SIM_RST, SIM_CLK);
    U74HC27 U19011(__A19_NET_240, CCH14, __A19_NET_241, GTONE, GOJAM, __A19_NET_242, GND, __A19_NET_248, __A19_NET_247, GTSET, GOJAM, __A19_NET_245, __A19_NET_248, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19012(__A19_NET_246, F5ASB2_n, __A19_NET_241, __A19_NET_247, __A19_NET_246, __A19_NET_248, GND, __A19_1__F5ASB0_n, __A19_NET_247, OTLNKM, __A19_NET_245, __A19_NET_248, __A19_NET_244, VCC, SIM_RST, SIM_CLK);
    U74HC02 U19013(CH1401, __A19_NET_244, RCH14_n, __A19_NET_232, __A19_NET_246, __A19_NET_235, GND, CA5_n, CXB7_n, __A19_NET_236, SB0_n, F05A_n, __A19_1__F5ASB0, VCC, SIM_RST, SIM_CLK);
    U74HC27 U19014(BR1_n, __A19_1__SH3MS_n, __A19_NET_234, __A19_1__SH3MS_n, BR1, __A19_1__OTLNK1, GND, __A19_NET_176, __A19_NET_238, __A19_1__UPL0_n, __A19_1__BLKUPL, __A19_NET_235, __A19_NET_234, VCC, SIM_RST, SIM_CLK);
    U74HC02 U19015(__A19_1__F5ASB2, F05A_n, SB2_n, __A19_1__F5BSB2, SB2_n, F05B_n, GND, __A19_1__XLNK0_n, __A19_NET_173, __A19_NET_172, __A19_1__XLNK1_n, __A19_NET_173, __A19_NET_171, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1) U19016(__A19_1__F5ASB2, F5ASB2_n, __A19_1__F5BSB2, F5BSB2_n, C45R, __A19_1__C45R_n, GND, __A19_NET_204, __A19_NET_162, __A19_NET_189, __A19_NET_207, __A19_1__UPL0_n, UPL0, VCC, SIM_RST, SIM_CLK);
    U74HC27 U19017(__A19_1__BLKUPL, __A19_NET_238, __A19_NET_168, __A19_NET_166, __A19_NET_182, INLNKM, GND, INLNKP, __A19_NET_167, __A19_NET_166, __A19_NET_182, __A19_NET_175, __A19_1__UPL1_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b0, 1'b0) U19018(__A19_NET_168, __A19_NET_176, __A19_NET_172, __A19_NET_167, __A19_NET_175, __A19_NET_171, GND, __A19_1__C45R_n, __A19_NET_181, __A19_NET_170, __A19_NET_170, __A19_NET_169, __A19_NET_181, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U19019(__A19_NET_178, __A19_NET_176, __A19_NET_175, __A19_NET_172, __A19_NET_171,  , GND,  , CA2_n, XB5_n, WOVR_n, OVF_n, T2P, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19020(__A19_NET_169, __A19_NET_170, __A19_NET_182, __A19_NET_182, __A19_NET_169, F04A, GND, BR1_n, __A19_1__C45R_n, __A19_1__UPRUPT, __A19_NET_169, __A19_NET_178, __A19_NET_179, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19021(__A19_NET_180, __A19_NET_179, __A19_NET_160, __A19_1__CH3311, __A19_NET_160, RCH33_n, GND, RCH33_n, __A19_1__BLKUPL, CH3310, CHWL05_n, WCH13_n, __A19_NET_158, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19022(__A19_NET_173, __A19_NET_158, __A19_NET_238, __A19_NET_238, __A19_NET_173, CCH13, GND, __A19_NET_173, CCH13, CH1305, WCH13_n, CHWL06_n, __A19_NET_159, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19023(__A19_NET_165, __A19_NET_159, __A19_NET_166, __A19_NET_166, __A19_NET_165, CCH13, GND, __A19_NET_165, CCH13, CH1306, CA5_n, XB5_n, __A19_NET_162, VCC, SIM_RST, SIM_CLK);
    U74HC27 U19024(__A19_NET_180, CCH33, CCHG_n, XT3_n, XB3_n, CCH33, GND, __A19_NET_164, __A19_NET_201, __A19_NET_203, CCH14, __A19_NET_160, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U19025(__A19_NET_196, __A19_NET_204, POUT_n, __A19_NET_199, __A19_NET_204, MOUT_n, GND, __A19_NET_204, ZOUT_n, __A19_NET_203, __A19_NET_163, __A19_NET_164, __A19_NET_201, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U19026(__A19_NET_163, WCH14_n, CHWL04_n, CH1404, RCH14_n, __A19_NET_201, GND, __A19_NET_201, F5ASB2_n, THRSTD, __A19_NET_196, __A19_NET_198, __A19_NET_197, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19027(__A19_NET_198, __A19_NET_197, __A19_NET_201, __A19_NET_202, __A19_NET_199, __A19_NET_200, GND, __A19_NET_202, __A19_NET_201, __A19_NET_200, __A19_NET_197, __A19_1__F5ASB0_n, __A19_1__THRSTp, VCC, SIM_RST, SIM_CLK);
    U74HC02 U19028(__A19_1__THRSTm, __A19_NET_202, __A19_1__F5ASB0_n, __A19_NET_207, CA5_n, XB6_n, GND, __A19_NET_189, POUT_n, __A19_NET_185, WCH14_n, CHWL05_n, __A19_NET_191, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U19029(__A19_NET_187, __A19_NET_189, MOUT_n, __A19_NET_190, __A19_NET_189, ZOUT_n, GND, __A19_NET_191, __A19_NET_205, __A19_NET_206, RCH14_n, __A19_NET_206, CH1405, VCC, SIM_RST, SIM_CLK);
    U74HC27 U19030(__A19_NET_206, __A19_NET_190, __A19_NET_255, __A19_NET_250, CCH14, __A19_NET_281, GND, __A19_NET_259, SB1_n, __A19_NET_297, __A19_NET_290, __A19_NET_205, CCH14, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U19031(EMSD, __A19_NET_206, F5ASB2_n, __A19_NET_184, __A19_NET_185, __A19_NET_186, GND, __A19_NET_184, __A19_NET_206, __A19_NET_186, __A19_NET_187, __A19_NET_188, __A19_NET_194, VCC, SIM_RST, SIM_CLK);
    U74HC02 U19032(__A19_NET_188, __A19_NET_194, __A19_NET_206, __A19_1__EMSp, __A19_NET_184, __A19_1__F5ASB0_n, GND, __A19_NET_194, __A19_1__F5ASB0_n, __A19_1__EMSm, CHWL09_n, WCH11_n, __A19_NET_326, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0) U19033(BLKUPL_n, __A19_1__BLKUPL, UPL1, __A19_1__UPL1_n, XLNK0, __A19_1__XLNK0_n, GND, __A19_1__XLNK1_n, XLNK1, __A19_2__OUTCOM, __A19_2__FF1109_n, __A19_2__ERRST, __A19_NET_285, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19034(__A19_2__FF1109_n, __A19_NET_326, __A19_NET_325, __A19_NET_325, __A19_2__FF1109_n, CCH11, GND, RCH11_n, __A19_2__FF1109_n, __A19_2__CH1109, CHWL10_n, WCH11_n, __A19_NET_286, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19035(__A19_2__FF1110_n, __A19_NET_286, __A19_NET_283, __A19_NET_283, __A19_2__FF1110_n, CCH11, GND, CAURST, __A19_NET_286, __A19_NET_285, RCH11_n, __A19_2__FF1110_n, __A19_2__CH1110, VCC, SIM_RST, SIM_CLK);
    U74HC04 U19036(__A19_2__FF1110_n, __A19_2__OT1110, __A19_2__FF1111_n, __A19_2__OT1111, __A19_2__FF1112_n, __A19_2__OT1112, GND, __A19_NET_262, __A19_NET_259, __A19_NET_261, __A19_NET_258, __A19_NET_260, __A19_NET_257, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19037(__A19_NET_280, CHWL11_n, WCH11_n, __A19_2__FF1111_n, __A19_NET_280, __A19_NET_284, GND, __A19_2__FF1111_n, CCH11, __A19_NET_284, RCH11_n, __A19_2__FF1111_n, __A19_2__CH1111, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19038(__A19_NET_279, CHWL12_n, WCH11_n, __A19_2__FF1112_n, __A19_NET_279, __A19_NET_278, GND, __A19_2__FF1112_n, CCH11, __A19_NET_278, RCH11_n, __A19_2__FF1112_n, __A19_2__CH1112, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19039(__A19_NET_282, CHWL10_n, WCH14_n, __A19_NET_255, __A19_NET_282, __A19_NET_281, GND, RCH14_n, __A19_NET_255, CH1410, CHWL09_n, WCH14_n, __A19_NET_293, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19040(__A19_NET_291, __A19_NET_293, __A19_NET_292, __A19_NET_292, __A19_NET_291, CCH14, GND, RCH14_n, __A19_NET_291, CH1409, CHWL08_n, WCH14_n, __A19_NET_298, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19041(__A19_NET_296, __A19_NET_298, __A19_NET_297, __A19_NET_297, __A19_NET_296, CCH14, GND, RCH14_n, __A19_NET_296, CH1408, CHWL07_n, WCH14_n, __A19_NET_295, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19042(__A19_NET_290, __A19_NET_295, __A19_NET_294, __A19_NET_294, __A19_NET_290, CCH14, GND, RCH14_n, __A19_NET_290, CH1407, CHWL06_n, WCH14_n, __A19_NET_287, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19043(__A19_NET_288, __A19_NET_287, __A19_NET_289, __A19_NET_289, __A19_NET_288, CCH14, GND, RCH14_n, __A19_NET_288, CH1406, __A19_NET_255, F5ASB2_n, GYROD, VCC, SIM_RST, SIM_CLK);
    U74HC27 U19044(SB1_n, __A19_NET_294, SB1_n, __A19_NET_296, __A19_NET_290, __A19_NET_257, GND, __A19_NET_253, __A19_NET_254, __A19_NET_249, __A19_NET_256, __A19_NET_258, __A19_NET_296, VCC, SIM_RST, SIM_CLK);
    U74HC02 U19045(__A19_2__GYENAB, SB1_n, __A19_NET_288, __A19_2__GYXP, __A19_NET_292, __A19_NET_262, GND, __A19_NET_262, __A19_NET_291, __A19_2__GYXM, __A19_NET_292, __A19_NET_261, __A19_2__GYYP, VCC, SIM_RST, SIM_CLK);
    U74HC02 U19046(__A19_2__GYYM, __A19_NET_261, __A19_NET_291, __A19_2__GYZP, __A19_NET_292, __A19_NET_260, GND, __A19_NET_260, __A19_NET_291, __A19_2__GYZM, CA4_n, XB7_n, __A19_NET_252, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0) U19047(__A19_NET_252, __A19_NET_251, __A19_NET_274, __A19_2__O44, F06B, __A19_2__F06B_n, GND, __A19_2__F07D_n, __A19_NET_268, __A19_2__F07C_n, __A19_NET_267, __A19_2__F7CSB1_n, __A19_NET_266, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U19048(__A19_NET_249, POUT_n, __A19_NET_251, __A19_NET_256, MOUT_n, __A19_NET_251, GND, ZOUT_n, __A19_NET_251, __A19_NET_250, __A19_NET_255, __A19_NET_253, __A19_NET_254, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U19049(__A19_2__GYRRST, F5ASB2_n, __A19_NET_254, __A19_2__GYRSET, F5ASB2_n, __A19_NET_253, GND, CHWL08_n, WCH13_n, __A19_NET_275, __A19_NET_275, __A19_NET_274, __A19_NET_273, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U19050(__A19_NET_274, __A19_NET_273, CCH13, CH1308, RCH13_n, __A19_NET_273, GND, WCH13_n, CHWL09_n, __A19_NET_272, __A19_NET_272, __A19_NET_277, __A19_NET_276, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19051(__A19_NET_269, __A19_NET_270, __A19_NET_311, CH1308, RCH13_n, __A19_NET_276, GND, __A19_NET_276, __A19_2__F07D_n, __A19_NET_265, FS07_n, __A19_2__F06B_n, __A19_NET_268, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U19052(__A19_NET_267, __A19_2__F06B_n, FS07A, __A19_NET_266, __A19_2__F07C_n, SB1_n, GND, __A19_NET_265, __A19_NET_264, __A19_NET_263, __A19_NET_263, F07B, __A19_NET_264, VCC, SIM_RST, SIM_CLK);
    U74HC27 U19053(SB2_n, __A19_NET_263, __A19_NET_276, CCH13, __A19_2__RHCGO, __A19_NET_277, GND, __A19_NET_318, __A19_NET_271, __A19_2__F07C_n, SB0_n, __A19_2__RHCGO, __A19_2__F07C_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0) U19054(__A19_NET_264, __A19_NET_271, SB2, __A19_2__CNTRSB_n, F10B, __A19_2__F10B_n, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U19055(SIGNX, __A19_2__F07C_n, SIGNY, __A19_2__F07C_n, __A19_2__F7CSB1_n, __A19_NET_322, GND, __A19_NET_320, SIGNZ, __A19_2__F07C_n, __A19_2__F7CSB1_n, __A19_NET_270, __A19_2__F7CSB1_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U19056(__A19_NET_311, __A19_NET_269, __A19_NET_318, __A19_NET_321, __A19_NET_322, __A19_NET_313, GND, __A19_NET_321, __A19_NET_318, __A19_NET_313, __A19_NET_320, __A19_NET_319, __A19_NET_317, VCC, SIM_RST, SIM_CLK);
    U74HC02 U19057(__A19_NET_319, __A19_NET_317, __A19_NET_318, __A19_NET_302, BMGXP, __A19_NET_315, GND, BMGXM, __A19_NET_312, __A19_NET_300, BMGYP, __A19_NET_316, __A19_NET_305, VCC, SIM_RST, SIM_CLK);
    U74HC27 U19058(F5ASB2_n, __A19_NET_269, F5ASB2_n, __A19_NET_311, GATEX_n, __A19_NET_312, GND, __A19_NET_316, F5ASB2_n, __A19_NET_321, GATEY_n, __A19_NET_315, GATEX_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U19059(F5ASB2_n, __A19_NET_313, F5ASB2_n, __A19_NET_317, GATEZ_n, __A19_NET_323, GND, __A19_NET_324, F5ASB2_n, __A19_NET_319, GATEZ_n, __A19_NET_314, GATEY_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 U19060(__A19_NET_303, BMGYM, __A19_NET_314, __A19_NET_304, BMGZP, __A19_NET_323, GND, BMGZM, __A19_NET_324, __A19_NET_299, __A19_2__O44, __A19_NET_302, BMAGXP, VCC, SIM_RST, SIM_CLK);
    U74HC02 U19061(BMAGXM, __A19_2__O44, __A19_NET_300, BMAGYP, __A19_2__O44, __A19_NET_305, GND, __A19_2__O44, __A19_NET_303, BMAGYM, __A19_2__O44, __A19_NET_304, BMAGZP, VCC, SIM_RST, SIM_CLK);
    U74HC02 U19062(BMAGZM, __A19_2__O44, __A19_NET_299, T1P, __A19_2__CNTRSB_n, __A19_2__F10B_n, GND, __A19_2__F10B_n, __A19_2__CNTRSB_n, T3P, F10A_n, __A19_2__CNTRSB_n, T5P, VCC, SIM_RST, SIM_CLK);
    U74HC27 U19063(FS10, F09B_n, __A19_2__F06B_n, T6ON_n, __A19_2__CNTRSB_n, T6P, GND,  ,  ,  ,  , T4P, __A19_2__CNTRSB_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20001(__A20_NET_148, CDUXP, __A20_NET_147, __A20_NET_147, __A20_NET_148, __A20_1__C1R, GND, CDUXM, __A20_NET_145, __A20_NET_150, __A20_NET_150, __A20_1__C1R, __A20_NET_145, VCC, SIM_RST, SIM_CLK);
    U74HC04 U20002(BKTF_n, __A20_NET_137, RSSB, __A20_NET_141, __A20_NET_170, __A20_1___CG2OUT, GND, __A20_1___CG5OUT, __A20_NET_162, __A20_NET_97, RSSB, __A20_NET_92, BKTF_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20003(__A20_NET_144, __A20_NET_147, __A20_NET_145, __A20_NET_146, __A20_NET_137, __A20_NET_144, GND, __A20_NET_146, __A20_NET_169, __A20_NET_151, __A20_NET_151, __A20_1__C1R, __A20_NET_169, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20004(C32A, __A20_1___CG1, __A20_NET_151, __A20_NET_140, CDUYP, __A20_NET_138, GND, __A20_NET_140, __A20_1__C2R, __A20_NET_138, CDUYM, __A20_NET_134, __A20_NET_139, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20005(__A20_NET_141, CA3_n, __A20_NET_148, CA3_n, CXB2_n, C32P, GND, C32M, __A20_NET_150, CA3_n, CXB2_n, __A20_1__C1R, CXB2_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20006(__A20_NET_134, __A20_NET_139, __A20_1__C2R, __A20_NET_135, __A20_NET_138, __A20_NET_134, GND, __A20_NET_137, __A20_NET_135, __A20_NET_136, __A20_NET_136, __A20_NET_168, __A20_NET_142, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U20007(__A20_NET_168, __A20_NET_142, __A20_1__C2R, __A20_NET_166, T2P, __A20_NET_167, GND, __A20_NET_166, __A20_1__C3R, __A20_NET_167, __A20_NET_137, __A20_NET_166, __A20_NET_176, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20008(__A20_NET_141, CA3_n, __A20_NET_140, CA3_n, CXB3_n, C33P, GND, C33M, __A20_NET_139, CA3_n, CXB3_n, __A20_1__C2R, CXB3_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20009(__A20_1___CG1, __A20_NET_169, __A20_1___CG1, __A20_NET_169, __A20_NET_168, __A20_NET_170, GND, __A20_1__C3R, __A20_NET_141, CA2_n, CXB4_n, C33A, __A20_NET_142, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U20010(__A20_NET_177, __A20_NET_176, __A20_NET_174, __A20_NET_174, __A20_NET_177, __A20_1__C3R, GND, GND, __A20_NET_177, C24A, T1P, __A20_NET_173, __A20_NET_172, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U20011(__A20_NET_173, __A20_NET_172, __A20_1__C4R, __A20_NET_156, __A20_NET_137, __A20_NET_172, GND, __A20_NET_156, __A20_NET_152, __A20_NET_157, __A20_NET_157, __A20_1__C4R, __A20_NET_152, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20012(__A20_NET_141, CA2_n, GND, __A20_NET_174, __A20_NET_157, C25A, GND, __A20_1__C5R, __A20_NET_141, CA2_n, CXB6_n, __A20_1__C4R, CXB5_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U20013(__A20_NET_154, T3P, __A20_NET_153, __A20_NET_153, __A20_NET_154, __A20_1__C5R, GND, __A20_NET_137, __A20_NET_154, __A20_NET_165, __A20_NET_165, __A20_NET_163, __A20_NET_164, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20014(__A20_NET_163, __A20_NET_164, __A20_1__C5R, __A20_NET_104, CDUZP, __A20_NET_103, GND, __A20_NET_104, __A20_1__C6R, __A20_NET_103, CDUZM, __A20_NET_101, __A20_NET_106, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U20015(C26A, GND, __A20_NET_174, __A20_NET_152, __A20_NET_164,  , GND,  , GND, __A20_NET_174, __A20_NET_152, __A20_NET_163, __A20_NET_162, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20016(__A20_NET_101, __A20_NET_106, __A20_1__C6R, __A20_NET_100, __A20_NET_103, __A20_NET_101, GND, __A20_NET_92, __A20_NET_100, __A20_NET_102, __A20_NET_102, __A20_NET_128, __A20_NET_107, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U20017(__A20_NET_128, __A20_NET_107, __A20_1__C6R, C34A, __A20_1___CG2OUT, __A20_NET_107, GND, TRNP, __A20_NET_94, __A20_NET_96, __A20_NET_96, __A20_1__C7R, __A20_NET_94, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20018(__A20_NET_97, CA3_n, __A20_NET_104, CA3_n, CXB4_n, C34P, GND, C34M, __A20_NET_106, CA3_n, CXB4_n, __A20_1__C6R, CXB4_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20019(__A20_NET_95, TRNM, __A20_NET_91, __A20_NET_91, __A20_NET_95, __A20_1__C7R, GND, __A20_NET_94, __A20_NET_91, __A20_NET_90, __A20_NET_92, __A20_NET_90, __A20_NET_93, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20020(__A20_NET_98, __A20_NET_93, __A20_NET_127, __A20_NET_127, __A20_NET_98, __A20_1__C7R, GND, T4P, __A20_NET_124, __A20_NET_122, __A20_NET_122, __A20_1__C8R, __A20_NET_124, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20021(__A20_NET_97, CA3_n, __A20_NET_96, CA3_n, CXB5_n, C35P, GND, C35M, __A20_NET_95, CA3_n, CXB5_n, __A20_1__C7R, CXB5_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20022(__A20_1___CG2OUT, __A20_NET_128, __A20_1___CG2OUT, __A20_NET_128, __A20_NET_127, __A20_NET_126, GND, __A20_1__C8R, __A20_NET_97, CA2_n, CXB7_n, C35A, __A20_NET_98, VCC, SIM_RST, SIM_CLK);
    U74HC04 U20023(__A20_NET_126, __A20_2___CG6, __A20_NET_118, __A20_1___CG1,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20024(__A20_NET_125, __A20_NET_92, __A20_NET_122, __A20_NET_133, __A20_NET_125, __A20_NET_132, GND, __A20_NET_133, __A20_1__C8R, __A20_NET_132, __A20_1___CG5OUT, __A20_NET_133, C27A, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U20025(__A20_NET_131, T5P, __A20_NET_129, __A20_NET_129, __A20_NET_131, __A20_1__C9R, GND, __A20_NET_92, __A20_NET_131, __A20_NET_111, __A20_NET_111, __A20_NET_115, __A20_NET_112, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U20026(__A20_NET_115, __A20_NET_112, __A20_1__C9R, __A20_NET_108, T6P, __A20_NET_109, GND, __A20_NET_108, __A20_1__C10R, __A20_NET_109, __A20_NET_92, __A20_NET_108, __A20_NET_121, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20027(__A20_NET_97, CA3_n, __A20_1___CG5OUT, __A20_NET_132, __A20_NET_112, C30A, GND, __A20_1__C10R, __A20_NET_97, CA3_n, CXB1_n, __A20_1__C9R, CXB0_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U20028(__A20_NET_119, __A20_NET_121, __A20_NET_120, __A20_NET_120, __A20_NET_119, __A20_1__C10R, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC4002 U20029(C31A, __A20_1___CG5OUT, __A20_NET_132, __A20_NET_115, __A20_NET_119,  , GND,  , __A20_1___CG5OUT, __A20_NET_132, __A20_NET_115, __A20_NET_120, __A20_NET_118, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20030(__A20_NET_236, PIPYP, __A20_NET_235, __A20_NET_235, __A20_NET_236, __A20_2__C1R, GND, PIPYM, __A20_NET_233, __A20_NET_238, __A20_NET_238, __A20_2__C1R, __A20_NET_233, VCC, SIM_RST, SIM_CLK);
    U74HC04 U20031(BKTF_n, __A20_NET_225, RSSB, __A20_NET_229, __A20_NET_259, CG13, GND, CG23, __A20_NET_250, __A20_NET_185, RSSB, __A20_NET_180, BKTF_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20032(__A20_NET_232, __A20_NET_235, __A20_NET_233, __A20_NET_234, __A20_NET_225, __A20_NET_232, GND, __A20_NET_234, __A20_NET_258, __A20_NET_239, __A20_NET_239, __A20_2__C1R, __A20_NET_258, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20033(C40A, __A20_2___CG1, __A20_NET_239, __A20_NET_228, PIPZP, __A20_NET_226, GND, __A20_NET_228, __A20_2__C2R, __A20_NET_226, PIPZM, __A20_NET_222, __A20_NET_227, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20034(__A20_NET_229, CA4_n, __A20_NET_236, CA4_n, CXB0_n, C40P, GND, C40M, __A20_NET_238, CA4_n, CXB0_n, __A20_2__C1R, CXB0_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20035(__A20_NET_222, __A20_NET_227, __A20_2__C2R, __A20_NET_223, __A20_NET_226, __A20_NET_222, GND, __A20_NET_225, __A20_NET_223, __A20_NET_224, __A20_NET_224, __A20_NET_257, __A20_NET_230, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U20036(__A20_NET_257, __A20_NET_230, __A20_2__C2R, __A20_NET_254, TRUND, __A20_NET_256, GND, __A20_NET_254, __A20_2__C3R, __A20_NET_256, __A20_NET_225, __A20_NET_254, __A20_NET_264, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20037(__A20_NET_229, CA4_n, __A20_NET_228, CA4_n, CXB1_n, C41P, GND, C41M, __A20_NET_227, CA4_n, CXB1_n, __A20_2__C2R, CXB1_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20038(__A20_2___CG1, __A20_NET_258, __A20_2___CG1, __A20_NET_258, __A20_NET_257, __A20_NET_259, GND, __A20_2__C3R, __A20_NET_229, CA5_n, CXB3_n, C41A, __A20_NET_230, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U20039(__A20_NET_265, __A20_NET_264, __A20_NET_263, __A20_NET_263, __A20_NET_265, __A20_2__C3R, GND, __A20_2___CG10OUT, __A20_NET_265, C53A, SHAFTD, __A20_NET_262, __A20_NET_261, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U20040(__A20_NET_262, __A20_NET_261, __A20_2__C4R, __A20_NET_243, __A20_NET_225, __A20_NET_261, GND, __A20_NET_243, __A20_NET_246, __A20_NET_244, __A20_NET_244, __A20_2__C4R, __A20_NET_246, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20041(__A20_NET_229, CA5_n, __A20_2___CG10OUT, __A20_NET_263, __A20_NET_244, C54A, GND, __A20_2__C5R, __A20_NET_229, CA5_n, CXB5_n, __A20_2__C4R, CXB4_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U20042(__A20_NET_241, THRSTD, __A20_NET_240, __A20_NET_240, __A20_NET_241, __A20_2__C5R, GND, __A20_NET_225, __A20_NET_241, __A20_NET_253, __A20_NET_253, __A20_NET_251, __A20_NET_252, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20043(__A20_NET_251, __A20_NET_252, __A20_2__C5R, __A20_NET_192, SHAFTP, __A20_NET_191, GND, __A20_NET_192, __A20_2__C6R, __A20_NET_191, SHAFTM, __A20_NET_189, __A20_NET_194, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U20044(C55A, __A20_2___CG10OUT, __A20_NET_263, __A20_NET_246, __A20_NET_252,  , GND,  , __A20_2___CG10OUT, __A20_NET_263, __A20_NET_246, __A20_NET_251, __A20_NET_250, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20045(__A20_NET_189, __A20_NET_194, __A20_2__C6R, __A20_NET_188, __A20_NET_191, __A20_NET_189, GND, __A20_NET_180, __A20_NET_188, __A20_NET_190, __A20_NET_190, __A20_NET_216, __A20_NET_195, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U20046(__A20_NET_216, __A20_NET_195, __A20_2__C6R, C36A, __A20_2___CG6, __A20_NET_195, GND, PIPXP, __A20_NET_182, __A20_NET_184, __A20_NET_184, __A20_2__C7R, __A20_NET_182, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20047(__A20_NET_185, CA3_n, __A20_NET_192, CA3_n, CXB6_n, C36P, GND, C36M, __A20_NET_194, CA3_n, CXB6_n, __A20_2__C6R, CXB6_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20048(__A20_NET_183, PIPXM, __A20_NET_179, __A20_NET_179, __A20_NET_183, __A20_2__C7R, GND, __A20_NET_182, __A20_NET_179, __A20_NET_178, __A20_NET_180, __A20_NET_178, __A20_NET_181, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20049(__A20_NET_186, __A20_NET_181, __A20_NET_215, __A20_NET_215, __A20_NET_186, __A20_2__C7R, GND, CDUXD, __A20_NET_212, __A20_NET_210, __A20_NET_210, __A20_2__C8R, __A20_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20050(__A20_NET_185, CA3_n, __A20_NET_184, CA3_n, CXB7_n, C37P, GND, C37M, __A20_NET_183, CA3_n, CXB7_n, __A20_2__C7R, CXB7_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20051(__A20_2___CG6, __A20_NET_216, __A20_2___CG6, __A20_NET_216, __A20_NET_215, __A20_NET_214, GND, __A20_2__C8R, __A20_NET_185, CA5_n, CXB0_n, C37A, __A20_NET_186, VCC, SIM_RST, SIM_CLK);
    U74HC04 U20052(__A20_NET_214, __A20_2___CG1, __A20_NET_206, __A20_2___CG10OUT,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20053(__A20_NET_213, __A20_NET_180, __A20_NET_210, __A20_NET_221, __A20_NET_213, __A20_NET_220, GND, __A20_NET_221, __A20_2__C8R, __A20_NET_220, CG26, __A20_NET_221, C50A, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U20054(__A20_NET_219, CDUYD, __A20_NET_217, __A20_NET_217, __A20_NET_219, __A20_2__C9R, GND, __A20_NET_180, __A20_NET_219, __A20_NET_199, __A20_NET_199, __A20_NET_203, __A20_NET_200, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U20055(__A20_NET_203, __A20_NET_200, __A20_2__C9R, __A20_NET_196, CDUZD, __A20_NET_197, GND, __A20_NET_196, __A20_2__C10R, __A20_NET_197, __A20_NET_180, __A20_NET_196, __A20_NET_209, VCC, SIM_RST, SIM_CLK);
    U74HC27 U20056(__A20_NET_185, CA5_n, CG26, __A20_NET_220, __A20_NET_200, C51A, GND, __A20_2__C10R, __A20_NET_185, CA5_n, CXB2_n, __A20_2__C9R, CXB1_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U20057(__A20_NET_207, __A20_NET_209, __A20_NET_208, __A20_NET_208, __A20_NET_207, __A20_2__C10R, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC4002 U20058(C52A, CG26, __A20_NET_220, __A20_NET_203, __A20_NET_207,  , GND,  , CG26, __A20_NET_220, __A20_NET_203, __A20_NET_208, __A20_NET_206, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21001(__A21_NET_204, C25A, C27A, C31A, C33A,  , GND,  , C35A, C37A, C41A, __A21_1__C43A, __A21_NET_203, VCC, SIM_RST, SIM_CLK);
    assign __A21_NET_205 = __A21_NET_205_U21002_2;
    assign __A21_NET_205 = __A21_NET_205_U21002_4;
    assign __A21_NET_205 = __A21_NET_205_U21002_6;
    assign __A21_NET_205 = __A21_NET_205_U21002_8;
    assign __A21_NET_147 = __A21_NET_147_U21002_10;
    assign __A21_NET_147 = __A21_NET_147_U21002_12;
    U74LVC07 U21002(__A21_NET_204, __A21_NET_205_U21002_2, __A21_NET_203, __A21_NET_205_U21002_4, __A21_NET_193, __A21_NET_205_U21002_6, GND, __A21_NET_205_U21002_8, __A21_NET_198, __A21_NET_147_U21002_10, __A21_NET_212, __A21_NET_147_U21002_12, __A21_NET_211, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21003(__A21_NET_193, __A21_1__C45A, __A21_1__C47A, C51A, C53A,  , GND,  , C26A, C27A, C32A, C33A, __A21_NET_212, VCC, SIM_RST, SIM_CLK);
    U74HC02 U21004(__A21_NET_198, C55A, __A21_1__C57A, __A21_NET_206, __A21_1__C56A, __A21_1__C57A, GND, __A21_1__30SUM, __A21_1__C60A, __A21_NET_222, __A21_1__50SUM, __A21_1__C60A, __A21_NET_220, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21005(__A21_NET_211, C36A, C37A, __A21_1__C42A, __A21_1__C43A,  , GND,  , __A21_1__C46A, __A21_1__C47A, C52A, C53A, __A21_NET_207, VCC, SIM_RST, SIM_CLK);
    assign __A21_NET_147 = __A21_NET_147_U21006_2;
    assign __A21_NET_147 = __A21_NET_147_U21006_4;
    assign __A21_NET_146 = __A21_NET_146_U21006_6;
    assign __A21_NET_146 = __A21_NET_146_U21006_8;
    assign __A21_NET_146 = __A21_NET_146_U21006_10;
    assign __A21_NET_146 = __A21_NET_146_U21006_12;
    U74LVC07 U21006(__A21_NET_207, __A21_NET_147_U21006_2, __A21_NET_206, __A21_NET_147_U21006_4, __A21_NET_209, __A21_NET_146_U21006_6, GND, __A21_NET_146_U21006_8, __A21_NET_172, __A21_NET_146_U21006_10, __A21_NET_173, __A21_NET_146_U21006_12, __A21_NET_168, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21007(__A21_NET_209, C24A, C25A, C26A, C27A,  , GND,  , C34A, C35A, C36A, C37A, __A21_NET_172, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21008(__A21_NET_173, __A21_1__C44A, __A21_1__C45A, __A21_1__C46A, __A21_1__C47A,  , GND,  , C54A, C55A, __A21_1__C56A, __A21_1__C57A, __A21_NET_168, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21009(__A21_NET_167, C30A, C31A, C32A, C33A,  , GND,  , C34A, C35A, C36A, C37A, __A21_NET_169, VCC, SIM_RST, SIM_CLK);
    assign __A21_1__32004K = __A21_1__32004K_U21010_2;
    assign __A21_1__32004K = __A21_1__32004K_U21010_4;
    assign __A21_NET_149 = __A21_NET_149_U21010_6;
    assign __A21_NET_149 = __A21_NET_149_U21010_8;
    assign __A21_NET_145 = __A21_NET_145_U21010_10;
    assign __A21_NET_145 = __A21_NET_145_U21010_12;
    U74LVC07 U21010(__A21_NET_167, __A21_1__32004K_U21010_2, __A21_NET_169, __A21_1__32004K_U21010_4, __A21_NET_189, __A21_NET_149_U21010_6, GND, __A21_NET_149_U21010_8, __A21_NET_183, __A21_NET_145_U21010_10, __A21_NET_182, __A21_NET_145_U21010_12, __A21_NET_222, VCC, SIM_RST, SIM_CLK);
    U74HC04 U21011(__A21_1__32004K, __A21_1__30SUM, __A21_NET_149, __A21_1__50SUM, DINC, DINC_n, GND, CXB0_n, XB0, CXB1_n, XB1, CXB2_n, XB2, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21012(__A21_NET_189, C50A, C51A, C52A, C53A,  , GND,  , C54A, C55A, __A21_1__C56A, __A21_1__C57A, __A21_NET_183, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21013(__A21_NET_182, C24A, C25A, C26A, C27A,  , GND,  , C40A, C41A, __A21_1__C42A, __A21_1__C43A, __A21_NET_184, VCC, SIM_RST, SIM_CLK);
    assign __A21_NET_223 = __A21_NET_223_U21015_2;
    assign __A21_NET_223 = __A21_NET_223_U21015_4;
    assign __A21_NET_223 = __A21_NET_223_U21015_6;
    assign __A21_NET_229 = __A21_NET_229_U21015_8;
    assign __A21_NET_229 = __A21_NET_229_U21015_10;
    assign __A21_NET_229 = __A21_NET_229_U21015_12;
    U74LVC07 U21015(__A21_NET_184, __A21_NET_223_U21015_2, __A21_NET_221, __A21_NET_223_U21015_4, __A21_NET_220, __A21_NET_223_U21015_6, GND, __A21_NET_229_U21015_8, __A21_NET_230, __A21_NET_229_U21015_10, __A21_NET_228, __A21_NET_229_U21015_12, __A21_NET_217, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21016(__A21_NET_221, __A21_1__C44A, __A21_1__C45A, __A21_1__C46A, __A21_1__C47A,  , GND,  , __A21_1__C45M, __A21_1__C46M, __A21_1__C57A, __A21_1__C60A, __A21_NET_153, VCC, SIM_RST, SIM_CLK);
    U74HC02 U21017(__A21_NET_148, __A21_1__30SUM, __A21_1__50SUM, CAD1, __A21_1__RSCT_n, __A21_NET_205, GND, __A21_1__RSCT_n, __A21_NET_147, CAD2, __A21_1__RSCT_n, __A21_NET_146, CAD3, VCC, SIM_RST, SIM_CLK);
    U74HC02 U21018(CAD4, __A21_1__RSCT_n, __A21_NET_148, CAD5, __A21_1__RSCT_n, __A21_NET_145, GND, __A21_1__RSCT_n, __A21_NET_223, CAD6, __A21_1__C45P, __A21_1__C46P, __A21_NET_152, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21019(C31A, __A21_1__C47A, C51A, C52A, C53A, __A21_NET_228, GND, __A21_NET_217, C54A, C55A, __A21_1__C56A, __A21_NET_230, C50A, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U21020(__A21_NET_155, INCSET_n, __A21_NET_153, __A21_NET_154, INCSET_n, __A21_NET_152, GND, INCSET_n, __A21_NET_229, __A21_NET_150, __A21_NET_155, __A21_1__SHINC, SHINC_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21021(__A21_1__SHINC, SHINC_n, T12A, SHANC_n, __A21_NET_154, __A21_1__SHANC, GND, SHANC_n, T12A, __A21_1__SHANC, __A21_NET_150, DINC, __A21_1__DINCNC_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U21022(DINC, __A21_1__DINCNC_n, T12A, __A21_NET_132, INCSET_n, __A21_NET_133, GND, __A21_NET_132, PINC, __A21_1__PINC_n, __A21_1__PINC_n, T12, PINC, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21023(__A21_NET_134, C24A, C25A, C26A, C27A,  , GND,  , C30A, C37P, C40P, C41P, __A21_NET_138, VCC, SIM_RST, SIM_CLK);
    assign __A21_NET_133 = __A21_NET_133_U21024_2;
    assign __A21_NET_133 = __A21_NET_133_U21024_4;
    assign __A21_NET_133 = __A21_NET_133_U21024_6;
    assign __A21_NET_142 = __A21_NET_142_U21024_8;
    assign __A21_NET_142 = __A21_NET_142_U21024_10;
    assign __A21_NET_157 = __A21_NET_157_U21024_12;
    U74LVC07 U21024(__A21_NET_134, __A21_NET_133_U21024_2, __A21_NET_138, __A21_NET_133_U21024_4, __A21_NET_144, __A21_NET_133_U21024_6, GND, __A21_NET_142_U21024_8, __A21_NET_141, __A21_NET_142_U21024_10, __A21_NET_140, __A21_NET_157_U21024_12, __A21_NET_161, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21025(__A21_1__C42P, __A21_1__C43P, __A21_1__C42M, __A21_1__C43M, __A21_1__C44M, __A21_NET_141, GND, __A21_NET_140, C37M, C40M, C41M, __A21_NET_144, __A21_1__C44P, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21026(__A21_NET_143, INCSET_n, __A21_NET_142, __A21_1__MINC_n, __A21_NET_143, MINC, GND, __A21_1__MINC_n, T12A, MINC, C35P, C36P, __A21_NET_158, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21027(C32P, C33P, C32M, C33M, C34M, __A21_NET_160, GND,  ,  ,  ,  , __A21_NET_161, C34P, VCC, SIM_RST, SIM_CLK);
    assign __A21_NET_157 = __A21_NET_157_U21028_2;
    assign __A21_NET_159 = __A21_NET_159_U21028_4;
    assign __A21_NET_159 = __A21_NET_159_U21028_6;
    U74LVC07 U21028(__A21_NET_158, __A21_NET_157_U21028_2, __A21_NET_160, __A21_NET_159_U21028_4, __A21_NET_164, __A21_NET_159_U21028_6, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21029(__A21_NET_162, INCSET_n, __A21_NET_157, __A21_1__PCDU_n, __A21_NET_162, PCDU, GND, __A21_1__PCDU_n, T12A, PCDU, C35M, C36M, __A21_NET_164, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21030(__A21_NET_163, INCSET_n, __A21_NET_159, __A21_1__MCDU_n, __A21_NET_163, MCDU, GND, __A21_1__MCDU_n, T12A, MCDU,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21031(__A21_NET_256, BMAGXP, __A21_NET_257, __A21_NET_257, __A21_NET_256, __A21_3__C42R, GND, BMAGXM, __A21_NET_263, __A21_NET_255, __A21_NET_255, __A21_3__C42R, __A21_NET_263, VCC, SIM_RST, SIM_CLK);
    U74HC04 U21032(BKTF_n, __A21_NET_242, RSSB, __A21_NET_243, __A21_NET_248, __A21_3__CG15, GND, CTROR, CTROR_n, __A21_NET_269, RSSB, __A21_NET_251, BKTF_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21033(__A21_NET_262, __A21_NET_257, __A21_NET_263, __A21_NET_258, __A21_NET_242, __A21_NET_262, GND, __A21_NET_258, __A21_NET_261, __A21_NET_259, __A21_NET_259, __A21_3__C42R, __A21_NET_261, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21034(__A21_1__C42A, CG13, __A21_NET_259, __A21_NET_238, BMAGYP, __A21_NET_239, GND, __A21_1__SHINC, __A21_1__SHANC, SHIFT_n, BMAGYM, __A21_NET_237, __A21_NET_235, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21035(__A21_NET_243, CA4_n, __A21_NET_256, CA4_n, CXB2_n, __A21_1__C42P, GND, __A21_1__C42M, __A21_NET_255, CA4_n, CXB2_n, __A21_3__C42R, CXB2_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21036(__A21_NET_237, __A21_NET_235, __A21_3__C43R, __A21_NET_234, __A21_NET_239, __A21_NET_237, GND, __A21_NET_242, __A21_NET_234, __A21_NET_231, __A21_NET_231, __A21_NET_233, __A21_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21037(__A21_NET_233, __A21_NET_232, __A21_3__C43R, __A21_NET_246, EMSD, __A21_NET_247, GND, __A21_NET_246, __A21_3__C56R, __A21_NET_247, __A21_NET_242, __A21_NET_246, __A21_NET_240, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21038(__A21_NET_243, CA4_n, __A21_NET_238, CA4_n, CXB3_n, __A21_1__C43P, GND, __A21_1__C43M, __A21_NET_235, CA4_n, CXB3_n, __A21_3__C43R, CXB3_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21039(CG13, __A21_NET_261, CG13, __A21_NET_261, __A21_NET_233, __A21_NET_248, GND, __A21_3__C56R, __A21_NET_243, CA5_n, CXB6_n, __A21_1__C43A, __A21_NET_232, VCC, SIM_RST, SIM_CLK);
    U74HC02 U2104( ,  ,  ,  ,  ,  , GND, __A21_NET_238, __A21_3__C43R, __A21_NET_239,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U21040(__A21_NET_241, __A21_NET_240, __A21_NET_276, __A21_NET_276, __A21_NET_241, __A21_3__C56R, GND, CG23, __A21_NET_241, __A21_1__C56A, OTLNKM, __A21_NET_245, __A21_NET_244, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U21041(__A21_NET_245, __A21_NET_244, __A21_3__C57R, __A21_NET_281, __A21_NET_242, __A21_NET_244, GND, __A21_NET_281, __A21_NET_277, __A21_NET_282, __A21_NET_282, __A21_3__C57R, __A21_NET_277, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21042(__A21_NET_243, CA5_n, CG23, __A21_NET_276, __A21_NET_282, __A21_1__C57A, GND, __A21_3__C60R, __A21_NET_243, CA6_n, CXB0_n, __A21_3__C57R, CXB7_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U21043(__A21_NET_286, ALTM, __A21_NET_280, __A21_NET_280, __A21_NET_286, __A21_3__C60R, GND, __A21_NET_242, __A21_NET_286, __A21_NET_283, __A21_NET_283, __A21_NET_285, __A21_NET_284, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21044(__A21_NET_285, __A21_NET_284, __A21_3__C60R, __A21_NET_300, BMAGZP, __A21_NET_279, GND, __A21_NET_300, __A21_3__C44R, __A21_NET_279, BMAGZM, __A21_NET_278, __A21_NET_299, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U21045(__A21_1__C60A, CG23, __A21_NET_276, __A21_NET_277, __A21_NET_284,  , GND,  , CG23, __A21_NET_276, __A21_NET_277, __A21_NET_285, CTROR_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21046(__A21_NET_278, __A21_NET_299, __A21_3__C44R, __A21_NET_298, __A21_NET_279, __A21_NET_278, GND, __A21_NET_251, __A21_NET_298, __A21_NET_296, __A21_NET_296, __A21_NET_297, __A21_NET_295, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U21047(__A21_NET_297, __A21_NET_295, __A21_3__C44R, __A21_1__C44A, __A21_3__CG15, __A21_NET_295, GND, INLNKP, __A21_NET_288, __A21_NET_287, __A21_NET_287, C45R, __A21_NET_288, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21048(__A21_NET_269, CA4_n, __A21_NET_300, CA4_n, CXB4_n, __A21_1__C44P, GND, __A21_1__C44M, __A21_NET_299, CA4_n, CXB4_n, __A21_3__C44R, CXB4_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21049(__A21_NET_294, INLNKM, __A21_NET_293, __A21_NET_293, __A21_NET_294, C45R, GND, __A21_NET_288, __A21_NET_293, __A21_NET_292, __A21_NET_251, __A21_NET_292, __A21_NET_289, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21050(__A21_NET_290, __A21_NET_289, __A21_NET_291, __A21_NET_291, __A21_NET_290, C45R, GND, RNRADP, __A21_NET_268, __A21_NET_253, __A21_NET_253, __A21_3__C46R, __A21_NET_268, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21051(__A21_NET_269, CA4_n, __A21_NET_287, CA4_n, CXB5_n, __A21_1__C45P, GND, __A21_1__C45M, __A21_NET_294, CA4_n, CXB5_n, C45R, CXB5_n, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21052(__A21_3__CG15, __A21_NET_297, __A21_3__CG15, __A21_NET_297, __A21_NET_291, __A21_NET_270, GND, __A21_3__C46R, __A21_NET_269, CA4_n, CXB6_n, __A21_1__C45A, __A21_NET_290, VCC, SIM_RST, SIM_CLK);
    U74HC04 U21053(__A21_NET_270, __A21_3__CG16, __A21_NET_266, CG26, XB3, CXB3_n, GND, CXB4_n, XB4, CXB5_n, XB5, CXB6_n, XB6, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21054(__A21_NET_272, __A21_NET_251, __A21_NET_273, __A21_NET_252, __A21_NET_272, __A21_NET_267, GND, __A21_NET_252, __A21_3__C46R, __A21_NET_267, __A21_3__CG16, __A21_NET_252, __A21_1__C46A, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21055(__A21_NET_254, RNRADM, __A21_NET_271, __A21_NET_271, __A21_NET_254, __A21_3__C46R, GND, __A21_NET_268, __A21_NET_271, __A21_NET_273,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21056( ,  ,  , __A21_NET_249, GYROD, __A21_NET_250, GND, __A21_NET_249, __A21_3__C47R, __A21_NET_250, __A21_NET_251, __A21_NET_249, __A21_NET_265, VCC, SIM_RST, SIM_CLK);
    U74HC27 U21057(__A21_NET_253, CA4_n, CA4_n, CXB6_n, __A21_NET_254, __A21_1__C46M, GND, __A21_3__C47R, __A21_NET_269, CA4_n, CXB7_n, __A21_1__C46P, CXB6_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U21058(__A21_NET_275, __A21_NET_265, __A21_NET_264, __A21_NET_264, __A21_NET_275, __A21_3__C47R, GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC27 U21059(__A21_3__CG16, __A21_NET_267, __A21_3__CG16, __A21_NET_267, __A21_NET_264, __A21_NET_266, GND,  ,  ,  ,  , __A21_1__C47A, __A21_NET_275, VCC, SIM_RST, SIM_CLK);
    U74HC04 U21060(XB7, CXB7_n, OCTAD2, CA2_n, OCTAD3, CA3_n, GND, CA4_n, OCTAD4, CA5_n, OCTAD5, CA6_n, OCTAD6, VCC, SIM_RST, SIM_CLK);
    U74HC04 U21061(SHIFT_n, SHIFT, RSCT, __A21_1__RSCT_n,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 U2062( ,  ,  ,  ,  ,  , GND, __A22_NET_194, CCH35, __A22_NET_193,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U22001(__A22_NET_125, __A22_1__DLKRPT, __A22_NET_124, DLKPLS, T10_n, __A22_NET_125, GND, __A22_NET_129, __A22_NET_122, __A22_1__DLKRPT, __A22_1__DLKRPT, __A22_NET_130, __A22_NET_122, VCC, SIM_RST, SIM_CLK);
    U74HC27 U22002(__A22_NET_125, DRPRST, __A22_NET_129, __A22_1__DLKRPT, __A22_NET_130, __A22_NET_128, GND, __A22_1__ADVCTR, __A22_1__RDOUT_n, __A22_1__WDORDR, __A22_1__BSYNC_n, __A22_NET_124, GOJAM, VCC, SIM_RST, SIM_CLK);
    U74HC04 U22003(DKEND, __A22_NET_129, __A22_NET_129, __A22_1__END, DKSTRT, __A22_NET_121, GND, __A22_1__DLKCLR, __A22_NET_121, __A22_NET_113, __A22_NET_111, __A22_1__DKCTR1_n, __A22_NET_118, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22004(__A22_NET_130, __A22_1__DLKRPT, __A22_NET_123, __A22_NET_123, __A22_NET_130, F10A, GND, __A22_NET_128, __A22_NET_127, __A22_NET_126, __A22_NET_126, CCH33, __A22_NET_127, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22005(CH3312, RCH33_n, __A22_NET_127, __A22_NET_111, __A22_1__DLKCLR, __A22_1__ADVCTR, GND, __A22_1__DLKCLR, __A22_NET_114, __A22_1__RDOUT_n, __A22_1__RDOUT_n, __A22_1__END, __A22_NET_114, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U22006(__A22_1__1CNT, __A22_NET_113, __A22_NET_109, __A22_NET_113, __A22_NET_116, __A22_NET_119, GND, __A22_NET_120, __A22_NET_118, __A22_1__DLKCLR, __A22_NET_119, __A22_NET_109, __A22_NET_119, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U22007(__A22_1__1CNT, __A22_NET_118, __A22_NET_109, __A22_NET_116, __A22_NET_119, __A22_NET_120, GND, __A22_NET_109, __A22_NET_120, __A22_NET_118, __A22_NET_141, __A22_NET_145, __A22_NET_117, VCC, SIM_RST, SIM_CLK);
    U74HC04 U22008(__A22_NET_120, __A22_1__DKCTR1, __A22_NET_141, __A22_1__DKCTR2_n, __A22_NET_142, __A22_1__DKCTR2, GND, __A22_1__DKCTR3_n, __A22_NET_148, __A22_1__DKCTR3, __A22_NET_146, __A22_1__DKCTR4_n, __A22_NET_134, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U22009(__A22_NET_117, __A22_NET_116, __A22_NET_145, __A22_NET_116, __A22_NET_144, __A22_NET_143, GND, __A22_NET_142, __A22_NET_141, __A22_1__DLKCLR, __A22_NET_143, __A22_NET_145, __A22_NET_143, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U22010(__A22_NET_144, __A22_NET_143, __A22_NET_142, __A22_NET_141, __A22_NET_145, __A22_NET_142, GND, __A22_NET_148, __A22_NET_150, __A22_NET_149, __A22_NET_151, __A22_NET_146, __A22_NET_147, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U22011(__A22_NET_149, __A22_NET_144, __A22_NET_150, __A22_NET_144, __A22_NET_147, __A22_NET_151, GND, __A22_NET_146, __A22_NET_148, __A22_1__DLKCLR, __A22_NET_151, __A22_NET_150, __A22_NET_151, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b0, 1'b1) U22012(__A22_NET_148, __A22_NET_150, __A22_NET_146, __A22_NET_133, __A22_NET_134, __A22_NET_139, GND, __A22_NET_140, __A22_NET_135, __A22_NET_132, __A22_NET_139, __A22_NET_135, __A22_NET_134, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U22013(__A22_NET_133, __A22_NET_147, __A22_NET_139, __A22_NET_147, __A22_NET_132, __A22_NET_140, GND, __A22_NET_135, __A22_NET_134, __A22_1__DLKCLR, __A22_NET_140, __A22_NET_139, __A22_NET_140, VCC, SIM_RST, SIM_CLK);
    U74HC04 U22014(__A22_NET_135, __A22_1__DKCTR4, __A22_NET_75, __A22_1__DKCTR5_n, __A22_NET_71, __A22_1__DKCTR5, GND, __A22_NET_83, __A22_1__BSYNC_n, __A22_NET_81, __A22_NET_80, __A22_NET_72, __A22_NET_81, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U22015(__A22_1__16CNT, __A22_NET_75, __A22_NET_137, __A22_1__32CNT, __A22_NET_138, __A22_NET_71, GND, __A22_NET_137, __A22_NET_71, __A22_NET_75, __A22_NET_83, __A22_NET_72, __A22_NET_62, VCC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U22016(__A22_1__16CNT, __A22_NET_132, __A22_NET_137, __A22_NET_132, __A22_1__32CNT, __A22_NET_138, GND, __A22_NET_71, __A22_NET_75, __A22_1__DLKCLR, __A22_NET_138, __A22_NET_137, __A22_NET_138, VCC, SIM_RST, SIM_CLK);
    U74HC02 U22017(__A22_NET_82, __A22_NET_62, __A22_NET_80, __A22_NET_80, __A22_NET_83, __A22_NET_82, GND, CHWL07_n, WCH13_n, __A22_NET_78, __A22_NET_77, __A22_NET_78, __A22_NET_79, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U22018(__A22_NET_77, CCH13, __A22_NET_79, CH1307, RCH13_n, __A22_NET_79, GND, __A22_1__DLKCLR, __A22_1__WDORDR, __A22_NET_63, __A22_NET_63, __A22_NET_62, __A22_1__WDORDR, VCC, SIM_RST, SIM_CLK);
    U74HC02 U22019(__A22_1__ORDRBT, __A22_NET_79, __A22_NET_63, __A22_NET_57, __A22_1__DKCTR5, __A22_1__DKCTR4, GND, __A22_1__DKCTR5, __A22_1__DKCTR4_n, __A22_NET_61, __A22_1__DKCTR4, __A22_1__DKCTR5_n, __A22_NET_58, VCC, SIM_RST, SIM_CLK);
    U74HC04 U22020(__A22_NET_57, __A22_1__HIGH0_n, __A22_NET_61, __A22_1__HIGH1_n, __A22_NET_58, __A22_1__HIGH2_n, GND, __A22_1__HIGH3_n, __A22_NET_69, __A22_1__LOW0_n, __A22_NET_65, __A22_1__LOW1_n, __A22_NET_66, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22021(__A22_NET_69, __A22_1__DKCTR4_n, __A22_1__DKCTR5_n, __A22_NET_103, CHWL16_n, WCH34_n, GND, __A22_NET_103, __A22_NET_102, __A22_NET_104, __A22_NET_104, CCH34, __A22_NET_102, VCC, SIM_RST, SIM_CLK);
    U74HC27 U22022(__A22_1__DKCTR1, __A22_1__DKCTR2, __A22_1__DKCTR1_n, __A22_1__DKCTR2, __A22_1__DKCTR3, __A22_NET_66, GND, __A22_NET_67, __A22_1__DKCTR1, __A22_1__DKCTR2_n, __A22_1__DKCTR3, __A22_NET_65, __A22_1__DKCTR3, VCC, SIM_RST, SIM_CLK);
    U74HC04 U22023(__A22_NET_67, __A22_1__LOW2_n, __A22_NET_101, __A22_1__LOW3_n, __A22_NET_97, __A22_1__LOW4_n, GND, __A22_1__LOW5_n, __A22_NET_98, __A22_1__LOW6_n, __A22_NET_107, __A22_1__LOW7_n, __A22_NET_108, VCC, SIM_RST, SIM_CLK);
    U74HC27 U22024(__A22_1__DKCTR1_n, __A22_1__DKCTR2_n, __A22_1__DKCTR1, __A22_1__DKCTR2, __A22_1__DKCTR3_n, __A22_NET_97, GND, __A22_NET_98, __A22_1__DKCTR1_n, __A22_1__DKCTR2, __A22_1__DKCTR3_n, __A22_NET_101, __A22_1__DKCTR3, VCC, SIM_RST, SIM_CLK);
    U74HC27 U22025(__A22_1__DKCTR1, __A22_1__DKCTR2_n, __A22_1__DKCTR1_n, __A22_1__DKCTR2_n, __A22_1__DKCTR3_n, __A22_NET_108, GND, __A22_NET_86, __A22_1__LOW0_n, __A22_NET_104, __A22_1__HIGH0_n, __A22_NET_107, __A22_1__DKCTR3_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22026(__A22_NET_90, WCH34_n, CHWL14_n, __A22_NET_88, __A22_NET_90, __A22_NET_89, GND, __A22_NET_88, CCH34, __A22_NET_89, __A22_1__DATA_n, __A22_1__WDORDR, __A22_NET_93, VCC, SIM_RST, SIM_CLK);
    U74HC27 U22027(__A22_1__HIGH0_n, __A22_NET_88, __A22_1__WRD1BP, __A22_1__WRD1B1, __A22_1__WRD2B2, __A22_NET_84, GND, __A22_NET_85, __A22_1__WRD2B3, __A22_NET_86, __A22_NET_87, __A22_NET_87, __A22_1__LOW1_n, VCC, SIM_RST, SIM_CLK);
    assign __A22_1__DATA_n = __A22_1__DATA_n_U22028_2;
    assign __A22_1__DATA_n = __A22_1__DATA_n_U22028_4;
    assign __A22_1__DATA_n = __A22_1__DATA_n_U22028_6;
    assign __A22_1__DATA_n = __A22_1__DATA_n_U22028_8;
    assign __A22_1__DATA_n = __A22_1__DATA_n_U22028_10;
    assign __A22_1__DATA_n = __A22_1__DATA_n_U22028_12;
    U74LVC07 U22028(__A22_NET_84, __A22_1__DATA_n_U22028_2, __A22_NET_85, __A22_1__DATA_n_U22028_4, __A22_NET_223, __A22_1__DATA_n_U22028_6, GND, __A22_1__DATA_n_U22028_8, __A22_NET_263, __A22_1__DATA_n_U22028_10, __A22_NET_249, __A22_1__DATA_n_U22028_12, __A22_NET_160, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22029(__A22_1__DKDAT_n, __A22_NET_93, __A22_1__ORDRBT, __A22_NET_234, WCH34_n, PC15_n, GND, __A22_NET_234, __A22_NET_235, __A22_NET_236, __A22_NET_236, CCH34, __A22_NET_235, VCC, SIM_RST, SIM_CLK);
    U74HC27 U22030(__A22_1__BSYNC_n, __A22_1__RDOUT_n, __A22_1__BSYNC_n, __A22_1__RDOUT_n, __A22_1__DKDAT_n, __A22_1__DKDATB, GND, __A22_1__WRD1BP, __A22_1__HIGH1_n, __A22_NET_236, __A22_1__LOW7_n, __A22_1__DKDATA, __A22_1__DKDAT_n, VCC, SIM_RST, SIM_CLK);
    U74HC04 U22031(DKBSNC, __A22_1__BSYNC_n,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22032(__A22_NET_232, WCH34_n, CHWL01_n, __A22_NET_231, __A22_NET_232, __A22_NET_233, GND, __A22_NET_231, CCH34, __A22_NET_233, WCH34_n, CHWL02_n, __A22_NET_242, VCC, SIM_RST, SIM_CLK);
    U74HC27 U22033(__A22_1__HIGH1_n, __A22_NET_231, __A22_1__HIGH1_n, __A22_NET_244, __A22_1__LOW5_n, __A22_NET_220, GND, __A22_NET_221, __A22_1__HIGH0_n, __A22_NET_239, __A22_1__LOW2_n, __A22_1__WRD1B1, __A22_1__LOW6_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U22034(__A22_NET_244, __A22_NET_242, __A22_NET_243, __A22_NET_243, __A22_NET_244, CCH34, GND, WCH34_n, CHWL13_n, __A22_NET_241, __A22_NET_241, __A22_NET_240, __A22_NET_239, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U22035(__A22_NET_223, __A22_NET_220, __A22_NET_221, __A22_NET_219, __A22_NET_230,  , GND,  , __A22_NET_264, __A22_NET_266, __A22_NET_268, __A22_NET_271, __A22_NET_263, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22036(__A22_NET_240, __A22_NET_239, CCH34, __A22_NET_222, WCH34_n, CHWL12_n, GND, __A22_NET_222, __A22_NET_216, __A22_NET_215, __A22_NET_215, CCH34, __A22_NET_216, VCC, SIM_RST, SIM_CLK);
    U74HC27 U22037(__A22_1__HIGH0_n, __A22_NET_215, __A22_1__HIGH0_n, __A22_NET_229, __A22_1__LOW4_n, __A22_NET_230, GND, __A22_NET_264, __A22_1__HIGH0_n, __A22_NET_224, __A22_1__LOW5_n, __A22_NET_219, __A22_1__LOW3_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22038(__A22_NET_217, WCH34_n, CHWL11_n, __A22_NET_229, __A22_NET_217, __A22_NET_218, GND, __A22_NET_229, CCH34, __A22_NET_218, WCH34_n, CHWL10_n, __A22_NET_228, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U22039(__A22_NET_224, __A22_NET_228, __A22_NET_225, __A22_NET_225, __A22_NET_224, CCH34, GND, WCH34_n, CHWL09_n, __A22_NET_227, __A22_NET_227, __A22_NET_226, __A22_NET_267, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22040(__A22_NET_226, __A22_NET_267, CCH34, __A22_NET_261, WCH34_n, CHWL08_n, GND, __A22_NET_261, __A22_NET_262, __A22_NET_265, __A22_NET_265, CCH34, __A22_NET_262, VCC, SIM_RST, SIM_CLK);
    U74HC27 U22041(__A22_1__HIGH0_n, __A22_NET_267, __A22_1__HIGH0_n, __A22_NET_265, __A22_1__LOW7_n, __A22_NET_268, GND, __A22_NET_271, __A22_1__HIGH1_n, __A22_NET_277, __A22_1__LOW0_n, __A22_NET_266, __A22_1__LOW6_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22042(__A22_NET_275, WCH34_n, CHWL07_n, __A22_NET_277, __A22_NET_275, __A22_NET_276, GND, __A22_NET_277, CCH34, __A22_NET_276, WCH34_n, CHWL06_n, __A22_NET_272, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U22043(__A22_NET_273, __A22_NET_272, __A22_NET_274, __A22_NET_274, __A22_NET_273, CCH34, GND, WCH34_n, CHWL05_n, __A22_NET_253, __A22_NET_253, __A22_NET_255, __A22_NET_254, VCC, SIM_RST, SIM_CLK);
    U74HC27 U22044(__A22_1__HIGH1_n, __A22_NET_273, __A22_1__HIGH1_n, __A22_NET_254, __A22_1__LOW2_n, __A22_NET_251, GND, __A22_NET_247, __A22_1__HIGH1_n, __A22_NET_260, __A22_1__LOW3_n, __A22_NET_248, __A22_1__LOW1_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22045(__A22_NET_255, __A22_NET_254, CCH34, __A22_NET_252, WCH34_n, CHWL04_n, GND, __A22_NET_252, __A22_NET_256, __A22_NET_260, __A22_NET_260, CCH34, __A22_NET_256, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U22046(__A22_NET_249, __A22_NET_248, __A22_NET_251, __A22_NET_247, __A22_NET_246,  , GND,  , __A22_NET_157, __A22_NET_158, __A22_NET_156, __A22_NET_168, __A22_NET_160, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22047(__A22_NET_259, WCH34_n, CHWL03_n, __A22_NET_257, __A22_NET_259, __A22_NET_258, GND, __A22_NET_257, CCH34, __A22_NET_258, WCH35_n, CHWL16_n, __A22_NET_172, VCC, SIM_RST, SIM_CLK);
    U74HC27 U22048(__A22_1__HIGH1_n, __A22_NET_257, __A22_1__HIGH2_n, __A22_NET_174, __A22_1__LOW0_n, __A22_NET_157, GND, __A22_NET_158, __A22_1__HIGH2_n, __A22_NET_171, __A22_1__LOW1_n, __A22_NET_246, __A22_1__LOW4_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U22049(__A22_NET_174, __A22_NET_172, __A22_NET_173, __A22_NET_173, __A22_NET_174, CCH35, GND, WCH35_n, CHWL14_n, __A22_NET_169, __A22_NET_169, __A22_NET_170, __A22_NET_171, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22050(__A22_NET_170, __A22_NET_171, CCH35, __A22_NET_180, WCH35_n, CHWL13_n, GND, __A22_NET_180, __A22_NET_181, __A22_NET_182, __A22_NET_182, CCH35, __A22_NET_181, VCC, SIM_RST, SIM_CLK);
    U74HC27 U22051(__A22_1__HIGH2_n, __A22_NET_182, __A22_1__HIGH2_n, __A22_NET_178, __A22_1__LOW3_n, __A22_NET_168, GND, __A22_NET_204, __A22_1__HIGH2_n, __A22_NET_152, __A22_1__LOW4_n, __A22_NET_156, __A22_1__LOW2_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22052(__A22_NET_176, WCH35_n, CHWL12_n, __A22_NET_178, __A22_NET_176, __A22_NET_179, GND, __A22_NET_178, CCH35, __A22_NET_179, WCH35_n, CHWL11_n, __A22_NET_159, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U22053(__A22_NET_152, __A22_NET_159, __A22_NET_153, __A22_NET_153, __A22_NET_152, CCH35, GND, WCH35_n, CHWL10_n, __A22_NET_154, __A22_NET_154, __A22_NET_155, __A22_NET_166, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22054(__A22_NET_155, __A22_NET_166, CCH35, __A22_NET_167, WCH35_n, CHWL09_n, GND, __A22_NET_167, __A22_NET_162, __A22_NET_161, __A22_NET_161, CCH35, __A22_NET_162, VCC, SIM_RST, SIM_CLK);
    U74HC27 U22055(__A22_1__HIGH2_n, __A22_NET_166, __A22_1__HIGH2_n, __A22_NET_161, __A22_1__LOW6_n, __A22_NET_208, GND, __A22_NET_207, __A22_1__HIGH2_n, __A22_NET_203, __A22_1__LOW7_n, __A22_NET_165, __A22_1__LOW5_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U22056(__A22_NET_201, __A22_NET_204, __A22_NET_165, __A22_NET_208, __A22_NET_207,  , GND,  , __A22_NET_187, __A22_NET_186, __A22_NET_185, __A22_NET_184, __A22_NET_183, VCC, SIM_RST, SIM_CLK);
    assign __A22_1__DATA_n = __A22_1__DATA_n_U22057_2;
    assign __A22_1__DATA_n = __A22_1__DATA_n_U22057_4;
    U74LVC07 U22057(__A22_NET_201, __A22_1__DATA_n_U22057_2, __A22_NET_183, __A22_1__DATA_n_U22057_4,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22058(__A22_NET_163, WCH35_n, CHWL08_n, __A22_NET_203, __A22_NET_163, __A22_NET_164, GND, __A22_NET_203, CCH35, __A22_NET_164, WCH35_n, CHWL07_n, __A22_NET_199, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U22059(__A22_NET_202, __A22_NET_199, __A22_NET_200, __A22_NET_200, __A22_NET_202, CCH35, GND, WCH35_n, CHWL06_n, __A22_NET_212, __A22_NET_212, __A22_NET_213, __A22_NET_214, VCC, SIM_RST, SIM_CLK);
    U74HC27 U22060(__A22_1__HIGH3_n, __A22_NET_202, __A22_1__HIGH3_n, __A22_NET_214, __A22_1__LOW1_n, __A22_NET_186, GND, __A22_NET_185, __A22_1__HIGH3_n, __A22_NET_211, __A22_1__LOW2_n, __A22_NET_187, __A22_1__LOW0_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22061(__A22_NET_213, __A22_NET_214, CCH35, __A22_NET_210, WCH35_n, CHWL05_n, GND, __A22_NET_210, __A22_NET_209, __A22_NET_211, __A22_NET_211, CCH35, __A22_NET_209, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22062(__A22_NET_192, WCH35_n, CHWL04_n, __A22_NET_194, __A22_NET_192, __A22_NET_193, GND,  ,  ,  , WCH35_n, CHWL03_n, __A22_NET_190, VCC, SIM_RST, SIM_CLK);
    U74HC27 U22063(__A22_1__HIGH3_n, __A22_NET_194, __A22_1__HIGH3_n, __A22_NET_198, __A22_1__LOW4_n, __A22_1__WRD2B3, GND, __A22_1__WRD2B2, __A22_1__HIGH3_n, __A22_NET_196, __A22_1__LOW5_n, __A22_NET_184, __A22_1__LOW3_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U22064(__A22_NET_198, __A22_NET_190, __A22_NET_191, __A22_NET_191, __A22_NET_198, CCH35, GND, WCH35_n, CHWL02_n, __A22_NET_197, __A22_NET_197, __A22_NET_195, __A22_NET_196, VCC, SIM_RST, SIM_CLK);
    U74HC02 U22065(__A22_NET_195, __A22_NET_196, CCH35,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
    assign SAP = SAP_U31001_29;
    assign SA08 = SA08_U31001_30;
    assign SA01 = SA01_U31001_31;
    assign SA09 = SA09_U31001_32;
    assign SA02 = SA02_U31001_33;
    assign SA10 = SA10_U31001_34;
    assign SA03 = SA03_U31001_35;
    assign SA11 = SA11_U31001_36;
    assign SA04 = SA04_U31001_38;
    assign SA12 = SA12_U31001_39;
    assign SA05 = SA05_U31001_40;
    assign SA13 = SA13_U31001_41;
    assign SA06 = SA06_U31001_42;
    assign SA14 = SA14_U31001_43;
    assign SA07 = SA07_U31001_44;
    assign SA16 = SA16_U31001_45;
    SST39VF200A U31001(__B01_1__FADDR16, __B01_1__FADDR15, __B01_1__FADDR14, __B01_1__FADDR13, __B01_1__FADDR12, __B01_1__FADDR11, __B01_1__FADDR10, __B01_1__FADDR9,  ,  , VCC,  ,  ,  ,  ,  ,  , __B01_1__FADDR8, __B01_1__FADDR7, __B01_1__FADDR6, __B01_1__FADDR5, __B01_1__FADDR4, __B01_1__FADDR3, __B01_1__FADDR2, __B01_1__FADDR1, __B01_NET_155, GND, __B01_NET_108, SAP_U31001_29, SA08_U31001_30, SA01_U31001_31, SA09_U31001_32, SA02_U31001_33, SA10_U31001_34, SA03_U31001_35, SA11_U31001_36, VCC, SA04_U31001_38, SA12_U31001_39, SA05_U31001_40, SA13_U31001_41, SA06_U31001_42, SA14_U31001_43, SA07_U31001_44, SA16_U31001_45, GND,  , GND, SIM_RST, SIM_CLK, EPCS_DATA, EPCS_CSN, EPCS_DCLK, EPCS_ASDI);
    U74HC04 U31002(ROPER, __B01_NET_181, ROPES, __B01_NET_182, ROPET, __B01_NET_144, GND, __B01_NET_171, STR14, __B01_NET_173, STR58, __B01_NET_142, STR912, VCC, SIM_RST, SIM_CLK);
    U74HC27 U31003(__B01_NET_144, LOMOD, ROPER, __B01_NET_141, __B01_NET_140, __B01_1__FADDR15, GND, __B01_NET_141, ROPES, LOMOD, STR14, __B01_1__FADDR16, STR14, VCC, SIM_RST, SIM_CLK);
    U74HC27 U31004(ROPET, HIMOD, ROPER, LOMOD, STR14, __B01_NET_149, GND, __B01_NET_148, ROPET, LOMOD, __B01_NET_171, __B01_NET_140, STR912, VCC, SIM_RST, SIM_CLK);
    U74HC02 U31005(__B01_NET_150, __B01_NET_182, __B01_NET_142, __B01_NET_147, __B01_NET_181, HIMOD, GND, HIMOD, STR58, __B01_NET_174, LOMOD, __B01_NET_173, __B01_NET_172, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U31006(__B01_1__FADDR14, __B01_NET_150, __B01_NET_149, __B01_NET_148, __B01_NET_147,  , GND,  , __B01_NET_177, __B01_NET_176, __B01_NET_180, __B01_NET_175, __B01_1__FADDR13, VCC, SIM_RST, SIM_CLK);
    U74HC27 U31007(ROPES, HIMOD, ROPES, LOMOD, STR14, __B01_NET_176, GND, __B01_NET_180, __B01_NET_182, HIMOD, __B01_NET_142, __B01_NET_177, STR912, VCC, SIM_RST, SIM_CLK);
    U74HC27 U31008(__B01_NET_182, LOMOD,  ,  ,  ,  , GND,  ,  ,  ,  , __B01_NET_175, __B01_NET_171, VCC, SIM_RST, SIM_CLK);
    U74HC02 U31009(__B01_1__FADDR12, __B01_NET_174, __B01_NET_172, __B01_1__FADDR11, STR210, STR19, GND, STR19, STR311, __B01_1__FADDR10, __B01_1__QUARTERB, __B01_1__QUARTERA, __B01_1__FADDR9, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31010(__B01_1__FADDR8, __B01_1__QUARTERA, __B01_1__QUARTERC, __B01_NET_99, __B01_NET_98, __B01_1__QUARTERA, GND, __B01_NET_99, __B01_1__CQA, __B01_1__QUARTERA, __B01_NET_92, __B01_NET_93, __B01_NET_98, VCC, SIM_RST, SIM_CLK);
    U74HC04 U31011(IL07, __B01_1__FADDR7, IL06, __B01_1__FADDR6, IL05, __B01_1__FADDR5, GND, __B01_1__FADDR4, IL04, __B01_1__FADDR3, IL03, __B01_1__FADDR2, IL02, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1) U31012(IL01, __B01_1__FADDR1, SBF, __B01_NET_108, SETAB, __B01_NET_92, GND, __B01_NET_93, RESETB, __B01_NET_223, __B01_NET_222, __B01_NET_104, __B01_NET_97, VCC, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U31013(__B01_NET_155, STR19, STR210, STR311, STR412,  , GND,  , XB1E, XB3E, XB5E, XB7E, __B01_2__ES01_n, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31014(__B01_NET_96, RESETA, __B01_NET_91, __B01_NET_94, __B01_NET_96, __B01_NET_97, GND, __B01_NET_94, RESETA, __B01_NET_97, __B01_NET_92, __B01_NET_130, __B01_NET_134, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1) U31015(__B01_NET_104, __B01_NET_105, __B01_NET_105, __B01_NET_106, __B01_NET_123, __B01_NET_102, GND, __B01_NET_103, __B01_NET_102, __B01_NET_101, __B01_NET_103, __B01_NET_121, __B01_NET_101, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1) U31016(__B01_NET_106, __B01_NET_91, RESETA, __B01_NET_130, SETCD, __B01_NET_139, GND, __B01_NET_138, RESETD, __B01_1__CQA, __B01_NET_137, __B01_NET_203, ZID, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U31017(__B01_NET_135, __B01_NET_134, __B01_1__QUARTERB, __B01_1__QUARTERB, __B01_NET_135, __B01_1__CQB, GND, __B01_NET_131, __B01_1__QUARTERC, __B01_NET_132, __B01_NET_132, __B01_1__CQC, __B01_1__QUARTERC, VCC, SIM_RST, SIM_CLK);
    U74HC02 U31018(__B01_NET_131, __B01_NET_139, __B01_NET_138, __B01_NET_137, CLROPE, __B01_NET_96, GND, YB1E, YB3E, __B01_2__ES07_n, YB2E, YB3E, __B01_2__ES08_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U31019(__B01_2__ES02_n, XB2E, XB3E, XB6E, XB7E,  , GND,  , XB4E, XB5E, XB6E, XB7E, __B01_2__ES03_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U31020(__B01_2__ES04_n, XT1E, XT3E, XT5E, XT7E,  , GND,  , XT2E, XT3E, XT6E, XT7E, __B01_2__ES05_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U31021(__B01_2__ES06_n, XT4E, XT5E, XT6E, XT7E,  , GND,  , YT1E, YT3E, YT5E, YT7E, __B01_2__ES09_n, VCC, SIM_RST, SIM_CLK);
    U74HC4002 U31022(__B01_2__ES10_n, YT2E, YT3E, YT6E, YT7E,  , GND,  , YT4E, YT5E, YT6E, YT7E, __B01_2__ES11_n, VCC, SIM_RST, SIM_CLK);
    assign SA07 = SA07_U31023_3;
    assign SA06 = SA06_U31023_5;
    assign SA05 = SA05_U31023_7;
    assign SA04 = SA04_U31023_9;
    assign SA03 = SA03_U31023_12;
    assign SA02 = SA02_U31023_14;
    assign SA01 = SA01_U31023_16;
    assign SAP = SAP_U31023_18;
    U74HC244 U31023(__B01_NET_203, GEMP, SA07_U31023_3, GEM01, SA06_U31023_5, GEM02, SA05_U31023_7, GEM03, SA04_U31023_9, GND, GEM04, SA03_U31023_12, GEM05, SA02_U31023_14, GEM06, SA01_U31023_16, GEM07, SAP_U31023_18, __B01_NET_203, VCC, SIM_RST, SIM_CLK);
    assign SA16 = SA16_U31024_3;
    assign SA14 = SA14_U31024_5;
    assign SA13 = SA13_U31024_7;
    assign SA12 = SA12_U31024_9;
    assign SA11 = SA11_U31024_12;
    assign SA10 = SA10_U31024_14;
    assign SA09 = SA09_U31024_16;
    assign SA08 = SA08_U31024_18;
    U74HC244 U31024(__B01_NET_203, GEM08, SA16_U31024_3, GEM09, SA14_U31024_5, GEM10, SA13_U31024_7, GEM11, SA12_U31024_9, GND, GEM12, SA11_U31024_12, GEM13, SA10_U31024_14, GEM14, SA09_U31024_16, GEM16, SA08_U31024_18, __B01_NET_203, VCC, SIM_RST, SIM_CLK);
    assign SAP = SAP_U31025_7;
    assign SA01 = SA01_U31025_8;
    assign SA02 = SA02_U31025_9;
    assign SA03 = SA03_U31025_10;
    assign SA04 = SA04_U31025_13;
    assign SA05 = SA05_U31025_14;
    assign SA06 = SA06_U31025_15;
    assign SA07 = SA07_U31025_16;
    assign SA08 = SA08_U31025_29;
    assign SA09 = SA09_U31025_30;
    assign SA10 = SA10_U31025_31;
    assign SA11 = SA11_U31025_32;
    assign SA12 = SA12_U31025_35;
    assign SA13 = SA13_U31025_36;
    assign SA14 = SA14_U31025_37;
    assign SA16 = SA16_U31025_38;
    MR0A16A U31025(__B01_2__RADDR1, __B01_2__RADDR2, __B01_2__RADDR3, __B01_2__RADDR4, __B01_2__RADDR5, GND, SAP_U31025_7, SA01_U31025_8, SA02_U31025_9, SA03_U31025_10, VCC, GND, SA04_U31025_13, SA05_U31025_14, SA06_U31025_15, SA07_U31025_16, __B01_NET_184, __B01_2__RADDR6, __B01_2__RADDR7, __B01_2__RADDR8, __B01_2__RADDR9, __B01_2__RADDR10, __B01_2__RADDR11, GND, GND, GND, VCC,  , SA08_U31025_29, SA09_U31025_30, SA10_U31025_31, SA11_U31025_32, VCC, GND, SA12_U31025_35, SA13_U31025_36, SA14_U31025_37, SA16_U31025_38, GND, GND, __B01_NET_187, GND, GND, GND, SIM_RST, SIM_CLK, SAP, SA01, SA02, SA03, SA04, SA05, SA06, SA07, SA08, SA09, SA10, SA11, SA12, SA13, SA14, SA16);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31026(__B01_NET_189, __B01_NET_185, __B01_NET_186, __B01_NET_235, __B01_2__ES01_n, __B01_NET_242, GND, __B01_NET_235, __B01_2__RADDR1, __B01_NET_188, __B01_NET_188, __B01_2__RESETK, __B01_2__RADDR1, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1) U31027(WEX, __B01_NET_185, WEY, __B01_NET_186, __B01_NET_189, __B01_NET_184, GND, __B01_NET_187, SBE, __B01_NET_242, SETEK, __B01_NET_220, __B01_NET_221, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31028(__B01_NET_238, __B01_2__ES02_n, __B01_NET_242, __B01_NET_237, __B01_NET_238, __B01_2__RADDR2, GND, __B01_NET_237, __B01_2__RESETK, __B01_2__RADDR2, __B01_2__ES03_n, __B01_NET_242, __B01_NET_240, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U31029(__B01_NET_239, __B01_NET_240, __B01_2__RADDR3, __B01_2__RADDR3, __B01_NET_239, __B01_2__RESETK, GND, __B01_2__ES04_n, __B01_NET_242, __B01_NET_224, __B01_NET_224, __B01_2__RADDR4, __B01_NET_227, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31030(__B01_2__RADDR4, __B01_NET_227, __B01_2__RESETK, __B01_NET_230, __B01_2__ES05_n, __B01_NET_242, GND, __B01_NET_230, __B01_2__RADDR5, __B01_NET_225, __B01_NET_225, __B01_2__RESETK, __B01_2__RADDR5, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31031(__B01_NET_233, __B01_2__ES06_n, __B01_NET_242, __B01_NET_232, __B01_NET_233, __B01_2__RADDR6, GND, __B01_NET_232, __B01_2__RESETK, __B01_2__RADDR6, __B01_2__ES07_n, __B01_NET_242, __B01_NET_244, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U31032(__B01_NET_243, __B01_NET_244, __B01_2__RADDR7, __B01_2__RADDR7, __B01_NET_243, __B01_2__RESETK, GND, __B01_2__ES08_n, __B01_NET_242, __B01_NET_198, __B01_NET_198, __B01_2__RADDR8, __B01_NET_197, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31033(__B01_2__RADDR8, __B01_NET_197, __B01_2__RESETK, __B01_NET_200, __B01_2__ES09_n, __B01_NET_242, GND, __B01_NET_200, __B01_2__RADDR9, __B01_NET_201, __B01_NET_201, __B01_2__RESETK, __B01_2__RADDR9, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31034(__B01_NET_190, __B01_2__ES10_n, __B01_NET_242, __B01_NET_192, __B01_NET_190, __B01_2__RADDR10, GND, __B01_NET_192, __B01_2__RESETK, __B01_2__RADDR10, __B01_2__ES11_n, __B01_NET_242, __B01_NET_204, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U31035(__B01_NET_205, __B01_NET_204, __B01_2__RADDR11, __B01_NET_116, CLROPE, __B01_NET_120, GND, __B01_NET_242, __B01_NET_219, __B01_2__RESETK, __B01_2__RESETK, __B01_NET_221, __B01_NET_214, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31036(__B01_NET_221, __B01_NET_214, __B01_NET_242, __B01_NET_120, RESETB, __B01_NET_121, GND, __B01_NET_120, __B01_NET_123, __B01_NET_119, __B01_NET_119, RESETB, __B01_NET_123, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1) U31037(__B01_NET_220, __B01_NET_222, __B01_NET_116, __B01_1__CQB, __B01_NET_223, __B01_NET_217, GND, __B01_NET_215, __B01_NET_217, __B01_NET_216, __B01_NET_215, __B01_NET_218, __B01_NET_216, VCC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1) U31038(__B01_NET_218, __B01_NET_219, __B01_NET_126, __B01_1__CQC, __B01_NET_124, __B01_NET_115, GND, __B01_NET_118, __B01_NET_115, __B01_NET_122, __B01_NET_118, __B01_NET_125, __B01_NET_122, VCC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31039(__B01_NET_126, CLROPE, __B01_NET_128, __B01_NET_128, RESETC, __B01_NET_125, GND, __B01_NET_128, __B01_NET_124, __B01_NET_129, __B01_NET_129, RESETC, __B01_NET_124, VCC, SIM_RST, SIM_CLK);
    U74HC02 U31040(__B01_2__RADDR11, __B01_NET_205, __B01_2__RESETK,  ,  ,  , GND,  ,  ,  ,  ,  ,  , VCC, SIM_RST, SIM_CLK);
endmodule
